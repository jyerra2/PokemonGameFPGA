module rand_gen();

endmodule

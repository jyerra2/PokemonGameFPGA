module user_pokeID(input logic [3:0] curr_level,
						 input logic [4:0] curr_ID,
						 output logic [4:0] new_ID);
//module gameState(   input Clk, Reset,
//						  input frameClk,
//						  input logic battle_done,
//						  input logic battle_start,
//						  
//						  
//						  
//						  output logic [1:0] curr_state
//						  
//						  
//						  
//						  );
//						  
//						  //battle_start from color mapper
//						  //battle_done from pokemon battle
//						  //curr_state(output of gameState) is used to indicate the state to the color mapper
//						  
//endmodule
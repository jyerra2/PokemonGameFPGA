//module Mem 2IO(  input logic Clk, 
//									 Reset,
//					 input logic [19:0] ADDR,
//					 input logic CE, UB, LB, OE, WE,
//					 input logic [15:0] selectMap,
//					 input logic [15:0] Data_from_SRAM,
//					 output logic [15:0] Data_to_ColorMapper,
//					 );
//					 
//					 
//					 always_comb
//					 begin
//					 Data_to_ColorMapper = Data_from_SRAM;
//					 end
//					 
//					 endmodule
//					 


//-------------------------------------------------------------------------
//    Color_Mapper.sv                                                    --
//    Stephen Kempf                                                      --
//    3-1-06                                                             --
//                                                                       --
//    Modified by David Kesler  07-16-2008                               --
//    Translated by Joe Meng    07-07-2013                               --
//    Modified by Po-Han Huang  03-03-2017                               --
//                                                                       --
//    Spring 2017 Distribution                                           --
//                                                                       --
//    For use with ECE 385 Lab 7                                         --
//    University of Illinois ECE Department                              --
//-------------------------------------------------------------------------


module  color_mapper (     input VGA_CLK, 
									Clk, frameClk,
                           input        [9:0] BallX, BallY,       // Ball coordinates

                           BallS,              // Ball size (defined in ball.sv)
                           DrawX, DrawY,
                           //input logic [2:0] gameControlBits,  //This is to select the background
                           input  logic [1:0] spriteDirControl,
                           input logic [3:0] counter,
                           // Coordinates of current drawing pixel
                           input [7:0] keycode,
                           input [15:0] Data,
				

                           output logic [2:0] pkmnChosen,

                           input logic [7:0] u [0:9],

                           input logic [7:0] w [0:9],

                           input logic [4:0] wildPokemonSprite,


                           input logic [5:0] hp_poke1,
                           hp_poke2,

                           output logic [1:0] curr_map,

                           input logic [3:0] battle_control,//from game_state which gets it from battle FSM

                           input logic [1:0] display_control,//from game_state

                           input logic [4:0] userPokemonSprite, //from userPkmnSelectModule

                           input logic [3:0] curr_level,//from Poke_Battle

                           output logic [4:0] PkmnChooseID, //This is to choose the ID of the Pokemon

                           output logic [7:0] VGA_R, VGA_G, VGA_B // VGA RGB output
                     );



logic ash_on;
logic [7:0] Red, Green, Blue;

//logic [2:0] pointer_on;

logic user_on;

//logic poke_select1, poke_select2, poke_select3;



/* The ball's (pixelated) circle is generated using the standard circle formula.  Note that while
   the single line is quite powerful descriptively, it causes the synthesis tool to use up three
   of the 12 available multipliers on the chip! Since the multiplicants are required to be signed,
   we have to first cast them from logic to int (signed by default) before they are multiplied. */

int DistX, DistY, Size;
assign DistX = DrawX - BallX;
assign DistY = DrawY - BallY;
//assign Size = BallS;

assign VGA_R = Red;
assign VGA_G = Green;
assign VGA_B = Blue;

//logic [7:0] MAP1[0:76799];
//logic [15:0] curr_map_pixel;


logic [7:0] ashDown0[0:1119];
logic [7:0] ashDown1[0:1119];
logic [7:0] ashDown2[0:1119];

logic [7:0] ashLeft0[0:1119];
logic [7:0] ashLeft1[0:1119];
logic [7:0] ashLeft2[0:1119];

logic [7:0] ashRight0[0:1119];
logic [7:0] ashRight1[0:1119];
logic [7:0] ashRight2[0:1119];

logic [7:0] ashUp0[0:1119];
logic [7:0] ashUp1[0:1119];
logic [7:0] ashUp2[0:1119];


logic [15:0] color;
logic [4:0] pokemon_id; //directly obtained from the color mapper
logic [7:0] spriteData;
logic [13:0] spriteAddr;

//
//logic [10:0] font_addr;
//logic [7:0] font_data;

logic [9:0] temp_X, temp_Y;
assign temp_X = DrawX;
assign temp_Y = DrawY;

logic [7:0] temp;

logic [4:0] pmknID;

always_ff
begin

//MAP1 = '{ 8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'hd,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h16,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h16,8'hd,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'h1,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h1,8'h1,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h1,8'hb,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'h1,8'hd,8'h4,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h14,8'hc,8'h1,8'hd,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'h14,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'h14,8'h14,8'hc,8'h1,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'h14,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h6,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'h1,8'h14,8'h14,8'hc,8'h1,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'h14,8'h13,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'ha,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h14,8'h14,8'hc,8'h1,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'h13,8'h14,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'hd,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'hd,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hd,8'hd,8'h13,8'h1,8'hd,8'h17,8'ha,8'ha,8'h17,8'h17,8'ha,8'ha,8'h17,8'h17,8'hd,8'h13,8'hd,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'hb,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hd,8'h1,8'h17,8'h17,8'ha,8'ha,8'h17,8'h17,8'hd,8'hd,8'h17,8'h17,8'h17,8'ha,8'h17,8'h17,8'h17,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'hb,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'h1,8'h17,8'ha,8'h17,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'h17,8'ha,8'h17,8'h16,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'hb,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'h16,8'ha,8'ha,8'h17,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h1,8'h17,8'ha,8'h1,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'h1,8'h17,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h1,8'h17,8'h1,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'h9,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h14,8'h14,8'h13,8'h1,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h16,8'h1,8'h4,8'h13,8'h14,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h14,8'h4,8'h13,8'h1,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h14,8'hc,8'hc,8'h4,8'h13,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h16,8'h1,8'h4,8'h14,8'h14,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h10,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h4,8'h13,8'hc,8'h13,8'h16,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hc,8'h9,8'h9,8'h9,8'h9,8'h9,8'h13,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h16,8'h4,8'h4,8'h14,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h1,8'h4,8'h4,8'h13,8'h14,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hc,8'h9,8'h4,8'h4,8'h13,8'h4,8'h9,8'h9,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h14,8'h14,8'h14,8'hc,8'h13,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h1,8'hd,8'h4,8'h4,8'h14,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h4,8'h4,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h14,8'h13,8'hc,8'hc,8'h13,8'h13,8'h14,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h4,8'h4,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h14,8'hc,8'h13,8'h1,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h1,8'h1,8'h1,8'h4,8'h4,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h14,8'hc,8'h9,8'h9,8'h4,8'h13,8'h13,8'h13,8'h13,8'h13,8'h1,8'h1,8'h13,8'h9,8'h9,8'h4,8'h1,8'h1,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h9,8'h9,8'h9,8'h14,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'hc,8'h13,8'h1,8'h1,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h1,8'h1,8'h1,8'hd,8'h14,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'hc,8'h9,8'hc,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h4,8'h4,8'h13,8'h4,8'h4,8'h13,8'h4,8'h4,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h4,8'h9,8'h9,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h13,8'h1,8'h1,8'h1,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h1,8'h1,8'h1,8'h1,8'hd,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h4,8'h9,8'h9,8'h4,8'h4,8'hc,8'h9,8'hc,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h1,8'h1,8'h1,8'h1,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h4,8'h9,8'h9,8'h9,8'h9,8'h4,8'hd,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'hd,8'h4,8'h4,8'hd,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h17,8'hd,8'hd,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hd,8'hd,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'hd,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'hd,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h1,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'hd,8'h10,8'ha,8'hd,8'h10,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'h4,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hd,8'h5,8'hd,8'h16,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hd,8'h5,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hc,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hc,8'hc,8'h4,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h1,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h16,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h4,8'hc,8'h9,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h10,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hc,8'hc,8'hc,8'h4,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h1,8'h16,8'h16,8'h16,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h16,8'h16,8'h16,8'h1,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hc,8'hc,8'h9,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hc,8'hc,8'hc,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'hd,8'ha,8'ha,8'hd,8'ha,8'h17,8'h17,8'h17,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h17,8'h17,8'h17,8'h17,8'hd,8'ha,8'ha,8'hd,8'h5,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'hc,8'hc,8'h9,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'h4,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hd,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'hc,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'ha,8'h4,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hd,8'ha,8'ha,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h4,8'hd,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'ha,8'ha,8'h4,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hd,8'ha,8'ha,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h10,8'ha,8'ha,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'hd,8'ha,8'ha,8'h4,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hd,8'ha,8'ha,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h5,8'ha,8'hd,8'hd,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'ha,8'hd,8'ha,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'hd,8'ha,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'ha,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'ha,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h4,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'ha,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'h7,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'h7,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'ha,8'ha,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h5,8'h5,8'h5,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'h5,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h7,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'h7,8'h5,8'h5,8'h5,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h5,8'h5,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'h5,8'h7,8'ha,8'ha,8'h11,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'ha,8'hf,8'ha,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h7,8'h5,8'hf,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'ha,8'h7,8'hf,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'ha,8'h11,8'ha,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h5,8'hf,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h7,8'h5,8'h7,8'hf,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'ha,8'ha,8'h11,8'h5,8'ha,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'h7,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'hf,8'ha,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'ha,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h11,8'ha,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'h17,8'hd,8'h4,8'h10,8'h5,8'h10,8'h5,8'h4,8'hd,8'h17,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'h7,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'h7,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'h7,8'hf,8'h11,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'h17,8'h17,8'h17,8'hd,8'h4,8'h7,8'h7,8'h7,8'h7,8'h5,8'hd,8'h17,8'h17,8'h17,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h11,8'ha,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'ha,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'h17,8'h17,8'h17,8'h17,8'h17,8'hd,8'h4,8'hd,8'h7,8'h7,8'h7,8'h10,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'h17,8'h17,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'hd,8'h1,8'hd,8'hd,8'hd,8'hd,8'h17,8'h17,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'h11,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'h17,8'h17,8'h17,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'h17,8'h17,8'h7,8'h7,8'h7,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h10,8'h10,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'ha,8'h7,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h7,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'ha,8'h10,8'h5,8'h5,8'h5,8'h10,8'ha,8'h7,8'h11,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'h7,8'hd,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h10,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h10,8'h10,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h10,8'h10,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h3,8'h5,8'h10,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h10,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h17,8'hd,8'hd,8'hd,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h1,8'h1,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h7,8'ha,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'ha,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'ha,8'hf,8'hf,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h10,8'h5,8'ha,8'h5,8'h7,8'hf,8'ha,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'h7,8'h7,8'hf,8'h7,8'h3,8'h5,8'h5,8'h5,8'h10,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h3,8'h17,8'h17,8'h17,8'h17,8'h3,8'ha,8'h11,8'ha,8'ha,8'h11,8'ha,8'ha,8'h11,8'ha,8'h3,8'h1,8'hd,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h17,8'h17,8'h17,8'h17,8'h1,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h1,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h17,8'h3,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h3,8'h17,8'h17,8'hd,8'h5,8'hd,8'h5,8'h5,8'hd,8'h5,8'hd,8'hd,8'h5,8'hd,8'h17,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h1,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'hd,8'hd,8'hd,8'hd,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'hd,8'h1,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h17,8'h7,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'hd,8'hd,8'hd,8'h5,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h10,8'hd,8'h17,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h17,8'h7,8'ha,8'he,8'he,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h17,8'h17,8'hd,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hd,8'h17,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'h7,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h1,8'h7,8'ha,8'h17,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'hd,8'hd,8'hd,8'h4,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h4,8'hd,8'hd,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h11,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'h11,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h1,8'hd,8'h17,8'h17,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'h17,8'h17,8'h1,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h17,8'h17,8'h17,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h17,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h7,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h7,8'h7,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'ha,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h7,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'h7,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h10,8'h5,8'h7,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h10,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'h7,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h10,8'h5,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'h7,8'hf,8'h11,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h11,8'ha,8'h10,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h7,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'h7,8'hf,8'h11,8'h7,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'ha,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h11,8'h11,8'ha,8'h7,8'ha,8'h10,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'h7,8'hf,8'ha,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h11,8'ha,8'h7,8'h7,8'h10,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'h11,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'ha,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'h11,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'ha,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'ha,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'ha,8'hf,8'hf,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hc,8'hc,8'h5,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h10,8'hc,8'hc,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h5,8'h8,8'hc,8'hc,8'h10,8'hd,8'ha,8'ha,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'ha,8'h5,8'hc,8'hc,8'h10,8'h8,8'hd,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h5,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h5,8'h7,8'hf,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h5,8'h5,8'hf,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'h5,8'hf,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h5,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h5,8'ha,8'hf,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'ha,8'h5,8'hf,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h5,8'hf,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h4,8'h4,8'hc,8'h10,8'hc,8'h10,8'ha,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'ha,8'ha,8'hc,8'hc,8'h10,8'h4,8'h4,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h7,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'h14,8'h4,8'h10,8'hc,8'h5,8'ha,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'h10,8'hc,8'h10,8'h4,8'h4,8'h10,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h4,8'h4,8'hc,8'h10,8'hc,8'h5,8'ha,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'hc,8'hc,8'h10,8'hc,8'h14,8'h4,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h12,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h14,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h14,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h14,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'ha,8'hf,8'h11,8'h7,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'h7,8'h7,8'h11,8'h7,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'ha,8'hf,8'h7,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'ha,8'hf,8'hf,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'h7,8'h7,8'h11,8'h7,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'h11,8'h7,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'ha,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h11,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h14,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'h7,8'h7,8'h10,8'h10,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'ha,8'h10,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h10,8'h10,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'h7,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h12,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'ha,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'ha,8'h10,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h10,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h10,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h14,8'h4,8'h10,8'h10,8'hc,8'h10,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h10,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'ha,8'h10,8'h10,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h10,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'hc,8'hc,8'h10,8'h8,8'h10,8'hc,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h4,8'h4,8'h4,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'hc,8'hc,8'h8,8'h8,8'hc,8'hc,8'hc,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hc,8'h4,8'h4,8'hc,8'h10,8'h8,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h9,8'h9,8'h9,8'h9,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h8,8'h8,8'hc,8'hc,8'h4,8'hc,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'h11,
//8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h4,8'h4,8'h4,8'hc,8'h10,8'h8,8'h8,8'h8,8'h8,8'h10,8'h9,8'h9,8'hc,8'hc,8'hc,8'h9,8'h9,8'h10,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'hc,8'h9,8'h4,8'h4,8'h4,8'h2,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h2,8'h5,8'hc,8'h4,8'h12,8'hc,8'hc,8'hc,8'hc,8'h10,8'h10,8'hc,8'h10,8'h10,8'hc,8'hc,8'h10,8'hc,8'h10,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'hc,8'hc,8'hc,8'hc,8'h4,8'h12,8'hc,8'hc,8'h8,8'h2,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'h11,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'h11,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'ha,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'h11,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h2,8'h8,8'hc,8'h4,8'h14,8'h14,8'h4,8'h9,8'h10,8'h2,8'h2,8'h2,8'hc,8'h9,8'hc,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h4,8'h9,8'h9,8'h4,8'h14,8'h12,8'hc,8'hc,8'h8,8'h2,8'h2,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h2,8'h8,8'h2,8'h8,8'h8,8'hc,8'h4,8'h4,8'h9,8'h9,8'h10,8'h5,8'hc,8'h10,8'h10,8'h9,8'h4,8'h10,8'hc,8'h10,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'hc,8'h9,8'hc,8'h4,8'h4,8'hc,8'h8,8'h8,8'h2,8'h8,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h2,8'h8,8'h2,8'h8,8'h5,8'h10,8'h10,8'h10,8'h10,8'h5,8'h10,8'h9,8'h9,8'hc,8'h10,8'hc,8'h9,8'h9,8'h4,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'h10,8'h10,8'h10,8'h10,8'h8,8'h8,8'h2,8'h8,8'h2,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'hc,8'h9,8'h9,8'h9,8'h9,8'h9,8'hc,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'hd,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'h5,8'h2,8'h8,8'h2,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h10,8'hc,8'hc,8'hc,8'h10,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h5,8'hd,8'hd,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'hd,8'h17,8'h5,8'h5,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h13,8'h17,8'h5,8'h5,8'hd,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hd,8'h5,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h2,8'h5,8'h5,8'hd,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h5,8'h7,8'hf,8'h7,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'h7,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'h5,8'hf,8'hf,8'h7,8'hf,8'h11,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'h7,8'hf,8'h7,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'h7,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'h7,8'hf,8'h7,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h13,8'hd,8'h17,8'hd,8'hd,8'hd,8'hd,8'h10,8'h5,8'h5,8'h5,8'hd,8'h12,8'h12,8'hd,8'h17,8'h17,8'hd,8'h13,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'hd,8'hd,8'h17,8'hd,8'h13,8'hd,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'ha,8'hd,8'h5,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'h10,8'hd,8'hd,8'hd,8'hd,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h10,8'h10,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h11,8'h7,8'h7,8'ha,8'h10,8'h5,8'h5,8'h10,8'h5,8'ha,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'h5,8'ha,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h11,8'h7,8'h7,8'h7,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'h17,8'h4,8'h4,8'h4,8'h17,8'h5,8'h10,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'h17,8'hd,8'h4,8'h4,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h17,8'h17,8'h17,8'hd,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'h5,8'ha,8'hd,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'ha,8'hc,8'h4,8'ha,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h10,8'h5,8'h5,8'ha,8'hf,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h10,8'h10,8'h5,8'ha,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'hd,8'h12,8'h13,8'hd,8'h17,8'ha,8'h10,8'h10,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h13,8'h12,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h4,8'h13,8'hd,8'h17,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'hc,8'h4,8'hd,8'h2,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h2,8'hd,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hc,8'h9,8'h4,8'ha,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h10,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'h11,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h10,8'ha,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h13,8'hd,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'h17,8'h13,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'hc,8'hc,8'h4,8'ha,8'h5,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hc,8'h9,8'h9,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'h4,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'h4,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'hc,8'hc,8'h4,8'ha,8'h2,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h2,8'ha,8'ha,8'ha,8'ha,8'hd,8'h10,8'h10,8'h10,8'h10,8'h10,8'h5,8'h4,8'hc,8'hc,8'h9,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h3,8'hd,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h17,8'h13,8'h4,8'hd,8'h17,8'h3,8'h17,8'h4,8'hd,8'h17,8'hd,8'h5,8'h5,8'hd,8'hd,8'h4,8'h13,8'h17,8'h17,8'h17,8'h4,8'h4,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hc,8'hc,8'hc,8'hd,8'ha,8'ha,8'hd,8'ha,8'ha,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'ha,8'ha,8'hd,8'h2,8'ha,8'hd,8'ha,8'ha,8'hd,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h5,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h17,8'h17,8'h4,8'h4,8'hd,8'h3,8'ha,8'h5,8'h5,8'hd,8'h17,8'hd,8'h17,8'h17,8'h3,8'hd,8'h4,8'hd,8'h17,8'h17,8'h5,8'h5,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'hd,8'h4,8'h13,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'h4,8'hc,8'hc,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h5,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h5,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'h11,8'h7,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'h7,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'h11,8'h7,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'ha,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h17,8'hd,8'hd,8'h17,8'hd,8'hd,8'h17,8'h3,8'hd,8'h5,8'h5,8'h5,8'h17,8'h3,8'hd,8'hd,8'h17,8'hd,8'hd,8'h17,8'h3,8'h17,8'h5,8'h5,8'h5,8'ha,8'h3,8'h17,8'h13,8'h17,8'hd,8'hd,8'h17,8'h3,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'ha,8'h4,8'hc,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h5,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h5,8'ha,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h11,8'hf,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h11,8'h11,8'h7,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h17,8'ha,8'hd,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h17,8'ha,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'ha,8'ha,8'hd,8'h17,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'ha,8'ha,8'h4,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h5,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h5,8'ha,8'ha,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'hd,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h5,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hd,8'ha,8'hd,8'hd,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'ha,8'hd,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'hd,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'hd,8'ha,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h13,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h13,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h13,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'ha,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'h12,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'hd,8'h17,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h10,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'h13,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h7,8'h5,8'ha,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'ha,8'h5,8'h5,8'h7,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h17,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h17,8'h13,8'h4,8'h13,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'h17,8'h5,8'h5,8'h5,8'h10,8'h5,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h10,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'h6,8'h7,8'h10,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h10,8'ha,8'h7,8'h7,8'h5,8'h10,8'h10,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h10,8'ha,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h10,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h10,8'h10,8'h5,8'h5,8'hd,8'hd,8'h17,8'h17,8'h13,8'h4,8'h12,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h10,8'h5,8'h17,8'hd,8'h17,8'h17,8'h4,8'h4,8'h13,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h17,8'hd,8'h17,8'h17,8'h4,8'h4,8'hd,8'h17,8'h5,8'h5,8'h10,8'h5,8'h5,8'hd,8'hd,8'h17,8'h17,8'h13,8'h4,8'h12,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'ha,8'h7,8'h6,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h7,8'h6,8'h6,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'hd,8'hd,8'hd,8'h17,8'h13,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h13,8'hd,8'h17,8'h3,8'h5,8'h10,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'hd,8'h13,8'hd,8'hd,8'h17,8'ha,8'h10,8'h10,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'h13,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h13,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h13,8'hd,8'h17,8'h3,8'h5,8'h5,8'h10,8'h10,8'hd,8'hd,8'hd,8'hd,8'hd,8'h13,8'hd,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'hd,8'h13,8'hd,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'h13,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h4,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h6,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h5,8'ha,8'h5,8'ha,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'h12,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h5,8'h10,8'h5,8'hd,8'h4,8'h4,8'h4,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'hd,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'h4,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'h4,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'hd,8'h13,8'h4,8'h4,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'hd,8'h5,8'h5,8'hd,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'ha,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'h4,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'ha,8'h5,8'h5,8'hd,8'hd,8'h4,8'h4,8'hd,8'h17,8'h3,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h3,8'hd,8'h12,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'h4,8'h17,8'h3,8'h17,8'h13,8'hd,8'h17,8'hd,8'h5,8'h5,8'hd,8'h13,8'h4,8'h4,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h3,8'hd,8'h13,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'h13,8'h17,8'h3,8'h17,8'h12,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h3,8'hd,8'h12,8'hd,8'h17,8'h5,8'h5,8'h5,8'h17,8'h4,8'h4,8'h4,8'h17,8'h17,8'h17,8'hd,8'hd,8'h17,8'hd,8'h5,8'h5,8'hd,8'hd,8'h4,8'h4,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h13,8'hd,8'h17,8'h3,8'hd,8'h4,8'h4,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h13,8'hd,8'h17,8'h17,8'h17,8'h4,8'h4,8'h17,8'h3,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h17,8'h17,8'h4,8'h4,8'hd,8'h3,8'hd,8'h5,8'h5,8'h17,8'hd,8'h13,8'h17,8'h17,8'h3,8'hd,8'h4,8'h13,8'h17,8'ha,8'h5,8'h5,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'hd,8'h4,8'h4,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h17,8'h17,8'h4,8'h4,8'hd,8'h3,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h17,8'h3,8'h4,8'h4,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h17,8'h17,8'h4,8'h4,8'hd,8'h3,8'hd,8'h5,8'h5,8'h17,8'hd,8'h13,8'h17,8'h17,8'h3,8'hd,8'h4,8'h13,8'h17,8'h17,8'h5,8'h5,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'hd,8'h4,8'h4,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'h13,8'h17,8'hd,8'h13,8'hd,8'h3,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'hd,8'h17,8'hd,8'h12,8'hd,8'h17,8'h3,8'h5,8'h5,8'h5,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'hd,8'h17,8'hd,8'h13,8'h17,8'h3,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'h13,8'h17,8'hd,8'h13,8'hd,8'h3,8'h17,8'h5,8'h5,8'h5,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'h5,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'hd,8'h17,8'hd,8'h13,8'h17,8'h3,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'h13,8'h17,8'hd,8'h13,8'hd,8'h3,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'hd,8'hd,8'h17,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h17,8'hd,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h7,8'h17,8'h7,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'hd,8'h17,8'h7,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'h7,8'h17,8'h7,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'h7,8'h17,8'h7,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h7,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'h7,8'h17,8'h7,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h7,8'h17,8'hd,8'h5,8'h5,8'hd,8'h17,8'h7,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h7,8'h17,8'h5,8'h5,8'h5,8'hd,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'h7,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'h7,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'ha,8'h5,8'hd,8'h13,8'h13,8'h7,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'ha,8'h5,8'hd,8'h12,8'hd,8'h7,8'h5,8'h17,8'h13,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'h5,8'ha,8'hd,8'h12,8'hd,8'h7,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'hd,8'h5,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'ha,8'h5,8'hd,8'h13,8'hd,8'h7,8'h5,8'h17,8'h13,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'h5,8'h5,8'hd,8'h12,8'hd,8'h7,8'h5,8'h17,8'h13,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'h5,8'ha,8'hd,8'h12,8'hd,8'h7,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'hd,8'h5,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h17,8'h5,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h3,8'h5,8'h5,8'h17,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'hd,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h17,8'h5,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h10,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h17,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h17,8'h5,8'h17,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h17,8'h5,8'h17,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h17,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h17,8'h5,8'h17,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h7,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h3,8'h3,8'h3,8'h3,8'hd,8'h17,8'h3,8'h3,8'h3,8'h7,8'ha,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'ha,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h7,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'ha,8'h3,8'h3,8'h3,8'h7,8'ha,8'h3,8'h3,8'h3,8'h3,8'hd,8'h3,8'h3,8'h3,8'h3,8'hd,8'h17,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h3,8'h3,8'h3,8'h3,8'hd,8'h7,8'h3,8'h3,8'h3,8'ha,8'ha,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'hd,8'hd,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h17,8'h3,8'h3,8'h3,8'hd,8'hd,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h3,8'h3,8'h3,8'h3,8'hd,8'h7,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'ha,8'h5,8'h7,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h3,8'ha,8'ha,8'ha,8'ha,8'h17,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h7,8'h17,8'h17,8'h17,8'h5,8'h5,8'hd,8'h17,8'h17,8'h17,8'hd,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h5,8'h17,8'hd,8'h13,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h10,8'hc,8'h9,8'h10,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'ha,8'hd,8'h13,8'hd,8'ha,8'h5,8'h5,8'h17,8'hd,8'h13,8'h17,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'ha,8'h3,8'hd,8'h3,8'ha,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'h5,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'ha,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h5,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h10,8'ha,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'ha,8'h3,8'hd,8'h3,8'ha,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'h5,8'ha,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'hd,8'h12,8'hd,8'h7,8'h5,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'h17,8'h13,8'h17,8'h7,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'ha,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'ha,8'h3,8'h17,8'h3,8'h7,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h17,8'h13,8'h17,8'ha,8'h10,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'ha,8'hd,8'h13,8'hd,8'h7,8'h5,8'h5,8'h17,8'hd,8'h12,8'h17,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'ha,8'h17,8'hd,8'h17,8'h3,8'h5,8'h5,8'h3,8'hd,8'hd,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'ha,8'h3,8'h3,8'h3,8'h7,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'ha,8'h17,8'h17,8'h17,8'ha,8'h10,8'h5,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'ha,8'hd,8'h13,8'hd,8'ha,8'h5,8'h5,8'h17,8'hd,8'h12,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'ha,8'h17,8'hd,8'h17,8'h7,8'h5,8'h5,8'h3,8'hd,8'hd,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'h3,8'h3,8'h3,8'h7,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'hd,8'h12,8'hd,8'h7,8'h5,8'h5,8'h3,8'hd,8'h13,8'h17,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'hd,8'h3,8'h7,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h10,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h10,8'hc,8'h9,8'h10,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'ha,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'ha,8'hd,8'hd,8'hd,8'h7,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'ha,8'h17,8'h13,8'h17,8'h3,8'h5,8'h5,8'h3,8'hd,8'hd,8'h3,8'ha,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'ha,8'h3,8'h17,8'h3,8'h7,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'ha,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'ha,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'h17,8'h12,8'h17,8'ha,8'h10,8'h5,8'h3,8'hd,8'h13,8'h17,8'ha,8'h5,8'ha,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'ha,8'h17,8'h12,8'h17,8'h7,8'h5,8'h5,8'h3,8'hd,8'h13,8'h3,8'ha,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'h17,8'h3,8'h7,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'h17,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h12,8'h17,8'ha,8'h5,8'h5,8'h3,8'hd,8'h12,8'h17,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h17,8'hd,8'h17,8'h7,8'h5,8'h5,8'h3,8'h17,8'hd,8'h3,8'ha,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'hc,8'h9,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'hd,8'hd,8'hd,8'hd,8'hd,8'h10,8'h5,8'hd,8'hd,8'hd,8'hd,8'h5,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'hc,8'h9};

// Main sprite/////ASH1 = '{ 8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h1,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h1,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h3,8'h3,8'h1,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h1,8'h1,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h3,8'h1,8'h1,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h1,8'h1,8'h1,8'h1,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h3,8'h1,8'h1,8'h1,8'h3,8'h7,8'h7,8'h7,8'h3,8'h2,8'h3,8'h7,8'h7,8'h7,8'h1,8'h1,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h3,8'h1,8'h1,8'h1,8'h3,8'h7,8'h3,8'h3,8'h2,8'h2,8'h3,8'h3,8'h7,8'h7,8'h1,8'h1,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h3,8'h1,8'h1,8'h1,8'h3,8'h7,8'h2,8'h3,8'h7,8'h7,8'h7,8'h2,8'h3,8'h7,8'h1,8'h1,8'h1,8'h3,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h1,8'h3,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h1,8'h1,8'h3,8'h3,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h1,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h3,8'h4,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h4,8'h4,8'h3,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h3,8'h5,8'h4,8'h4,8'h5,8'h4,8'h7,8'h3,8'h5,8'h5,8'h4,8'h7,8'h4,8'h5,8'h4,8'h4,8'h4,8'h4,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h3,8'h4,8'h4,8'h4,8'h5,8'h4,8'h7,8'h3,8'h5,8'h5,8'h4,8'h7,8'h3,8'h5,8'h4,8'h4,8'h4,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h3,8'h3,8'h4,8'h4,8'h4,8'h3,8'h4,8'h5,8'h5,8'h4,8'h3,8'h4,8'h4,8'h4,8'h4,8'h4,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h3,8'h3,8'h4,8'h1,8'h4,8'h5,8'h5,8'h4,8'h1,8'h4,8'h4,8'h3,8'h3,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h1,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h1,8'h4,8'h3,8'h7,8'h7,8'h7,8'h3,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h4,8'h4,8'h3,8'h0,8'h0,8'h0,8'h0,8'h3,8'h4,8'h5,8'h3,8'h7,8'h7,8'h7,8'h3,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h3,8'h7,8'h7,8'h3,8'h5,8'h4,8'h3,8'h0,8'h0,8'h0,8'h0,8'h3,8'h1,8'h5,8'h4,8'h4,8'h3,8'h7,8'h3,8'h6,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h6,8'h6,8'h3,8'h7,8'h3,8'h4,8'h5,8'h4,8'h3,8'h0,8'h0,8'h0,8'h0,8'h3,8'h1,8'h1,8'h4,8'h4,8'h3,8'h7,8'h3,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h7,8'h7,8'h3,8'h4,8'h4,8'h1,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h6,8'h6,8'h3,8'h1,8'h1,8'h3,8'h6,8'h6,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h0,8'h0,8'h0,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h7,8'h7,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0};
//ASH1 = '{8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h1,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h1,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h16,8'h16,8'h1,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h1,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h1,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'hb,8'hb,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'h11,8'h3,8'h3,8'h3,8'h3,8'h9,8'h11,8'h11,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h11,8'h11,8'h9,8'h3,8'h3,8'h3,8'h3,8'h11,8'hb,8'hb,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'h3,8'hb,8'hb,8'hb,8'hb,8'h9,8'h11,8'h11,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h11,8'h11,8'h9,8'h3,8'h3,8'hb,8'hb,8'h3,8'hb,8'hb,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h9,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'h9,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h9,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'h9,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h1,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h1,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h3,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h17,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h3,8'hd,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'hd,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h4,8'h9,8'h4,8'h3,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h7,8'h9,8'h9,8'h4,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'hd,8'h9,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h3,8'h9,8'hd,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h4,8'h4,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h3,8'h11,8'h9,8'hd,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h7,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'hd,8'h3,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h9,8'h9,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'h11,8'h3,8'h11,8'h11,8'h9,8'h9,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h9,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h2,8'h2,8'h11,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'h2,8'h11,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h9,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h9,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h9,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h9,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h9,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h9,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h9,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hb,8'hb,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hf,8'hf,8'hf,8'hf,8'h11,8'h3,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h11,8'h11,8'h11,8'h11,8'h11,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h11,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hf,8'hf,8'hf,8'h11,8'h7,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h11,8'hf,8'hf,8'hf,8'hf,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'hf,8'hf,8'h11,8'h17,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h3,8'h11,8'hf,8'hf,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h17,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h3,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h0,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h0,8'h0,8'h0,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h11,8'h11,8'h16,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h11,8'h11,8'h16,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h16,8'h3,8'h3,8'h16,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h16,8'h3,8'h3,8'h16,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0};

ashDown0 = '{ 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h1, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h15, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h11, 8'h16, 8'h16, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h1, 8'h16, 8'h11, 8'h11, 8'h15, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h11, 8'h16, 8'h1, 8'h3, 8'h11, 8'h11, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'h13, 8'hd, 8'hd, 8'h11, 8'hd, 8'hd, 8'hd, 8'h11, 8'hd, 8'hd, 8'h13, 8'h17, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h13, 8'h13, 8'h14, 8'h14, 8'h3, 8'h14, 8'h14, 8'h14, 8'h3, 8'h14, 8'h14, 8'h13, 8'h13, 8'hd, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h13, 8'h17, 8'h14, 8'h14, 8'h14, 8'h17, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'hd, 8'h13, 8'h13, 8'h17, 8'h14, 8'h14, 8'h14, 8'h17, 8'h13, 8'h13, 8'hd, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h17, 8'h11, 8'h11, 8'h2, 8'h2, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h2, 8'h2, 8'h11, 8'h11, 8'h11, 8'hd, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h14, 8'h13, 8'h17, 8'h11, 8'h2, 8'h2, 8'ha, 8'ha, 8'ha, 8'ha, 8'ha, 8'h2, 8'h2, 8'h11, 8'h17, 8'hd, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h14, 8'h11, 8'h2, 8'h2, 8'h8, 8'h8, 8'h8, 8'h8, 8'h8, 8'h2, 8'h2, 8'h11, 8'h14, 8'h14, 8'h13, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'hd, 8'h11, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h11, 8'hd, 8'hd, 8'h13, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h11, 8'h11, 8'h2, 8'h2, 8'h2, 8'h16, 8'h16, 8'h16, 8'h2, 8'h2, 8'h2, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
           ashDown1 = ' { 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h1, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h15, 8'h15, 8'h7, 8'h11, 8'h11, 8'h3, 8'h16, 8'h1, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h15, 8'h15, 8'h7, 8'h11, 8'h11, 8'h3, 8'h16, 8'h1, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h1, 8'h16, 8'h3, 8'h11, 8'h15, 8'h11, 8'h11, 8'h7, 8'h15, 8'h11, 8'h3, 8'h16, 8'h1, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h13, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h13, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h13, 8'h13, 8'h14, 8'h14, 8'h3, 8'h14, 8'h14, 8'h17, 8'h3, 8'h14, 8'h13, 8'h13, 8'hd, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h13, 8'h13, 8'h14, 8'h14, 8'h3, 8'h14, 8'h14, 8'h17, 8'h3, 8'h14, 8'h13, 8'h13, 8'hd, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h13, 8'h13, 8'h17, 8'h14, 8'h14, 8'hd, 8'h17, 8'h13, 8'h13, 8'h13, 8'h17, 8'h11, 8'h17, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h13, 8'h13, 8'h17, 8'h14, 8'h14, 8'hd, 8'h17, 8'h13, 8'h13, 8'h13, 8'h17, 8'h11, 8'h17, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'hd, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h17, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'ha, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'ha, 8'h2, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'ha, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'ha, 8'h2, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h14, 8'h14, 8'hd, 8'h17, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h13, 8'h13, 8'h1, 8'h17, 8'h2, 8'h16, 8'h16, 8'h16, 8'h2, 8'h8, 8'ha, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h13, 8'h13, 8'h1, 8'h17, 8'h2, 8'h16, 8'h16, 8'h16, 8'h2, 8'h8, 8'ha, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
ashDown2 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h16, 8'h16, 8'h11, 8'h11, 8'h7, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'hd, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h3, 8'h13, 8'h13, 8'h14, 8'hd, 8'h3, 8'h14, 8'h14, 8'h12, 8'h11, 8'h14, 8'h13, 8'h13, 8'h13, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h3, 8'h13, 8'h13, 8'h14, 8'hd, 8'h3, 8'h14, 8'h14, 8'h12, 8'h11, 8'h14, 8'h13, 8'h13, 8'h13, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h17, 8'h11, 8'h17, 8'hd, 8'h13, 8'hd, 8'hd, 8'h14, 8'h14, 8'h14, 8'h17, 8'h13, 8'h13, 8'h1, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h17, 8'h11, 8'h17, 8'hd, 8'h13, 8'hd, 8'hd, 8'h14, 8'h14, 8'h14, 8'h17, 8'h13, 8'h13, 8'h1, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h17, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h2, 8'h8, 8'ha, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h2, 8'h8, 8'ha, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h3, 8'hd, 8'h14, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h2, 8'h2, 8'hd, 8'h16, 8'h16, 8'h16, 8'h2, 8'h17, 8'hd, 8'h13, 8'h13, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h2, 8'h2, 8'hd, 8'h16, 8'h16, 8'h16, 8'h2, 8'h17, 8'hd, 8'h13, 8'h13, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0 };

           ashLeft0 = ' {8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h15, 8'h15, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h1, 8'h1, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h3, 8'h3, 8'h17, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h1, 8'h17, 8'h17, 8'h17, 8'h1, 8'h17, 8'h17, 8'h17, 8'h1, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h11, 8'h13, 8'h13, 8'h13, 8'h17, 8'h14, 8'h13, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h11, 8'h13, 8'h13, 8'h13, 8'h17, 8'h14, 8'h13, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h14, 8'h14, 8'h3, 8'h14, 8'h13, 8'h13, 8'hd, 8'h14, 8'h13, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'hd, 8'h14, 8'h13, 8'h13, 8'h14, 8'h13, 8'hd, 8'hd, 8'h7, 8'h11, 8'h11, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'hd, 8'hd, 8'hd, 8'hd, 8'h17, 8'h3, 8'h17, 8'h17, 8'h15, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h17, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h8, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'ha, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'hd, 8'h7, 8'h7, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h14, 8'h14, 8'h14, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'hd, 8'hd, 8'hd, 8'h11, 8'h11, 8'h11, 8'h7, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h3, 8'h3, 8'h3, 8'h17, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
ashLeft1 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h15, 8'h7, 8'h11, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h15, 8'h7, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h15, 8'h7, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h17, 8'h1, 8'h1, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h3, 8'h3, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h1, 8'h3, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h14, 8'h3, 8'h17, 8'h14, 8'h13, 8'h17, 8'h14, 8'h14, 8'h14, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h17, 8'h14, 8'h17, 8'hd, 8'h14, 8'h13, 8'h13, 8'h14, 8'h14, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'hd, 8'h13, 8'h13, 8'h13, 8'h13, 8'hd, 8'hd, 8'h1, 8'h7, 8'h7, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h17, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'hd, 8'hd, 8'hd, 8'h17, 8'h17, 8'h17, 8'h17, 8'hd, 8'h15, 8'h15, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h17, 8'h17, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h13, 8'h12, 8'h13, 8'h11, 8'h11, 8'h11, 8'h2, 8'h2, 8'h15, 8'h15, 8'h15, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h11, 8'h14, 8'h14, 8'h12, 8'h11, 8'h11, 8'h11, 8'h2, 8'h8, 8'h15, 8'h15, 8'he, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h14, 8'h14, 8'h13, 8'h11, 8'h11, 8'h11, 8'h2, 8'h2, 8'h7, 8'h17, 8'he, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h13, 8'h13, 8'hd, 8'h11, 8'h11, 8'h11, 8'h2, 8'h2, 8'h11, 8'h17, 8'he, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
           ashLeft2 = ' {8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h17, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h1, 8'h15, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h1, 8'h15, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h17, 8'h3, 8'h3, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h1, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h1, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h16, 8'h3, 8'h3, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h3, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h17, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h17, 8'h17, 8'h11, 8'h3, 8'h17, 8'h17, 8'h3, 8'h3, 8'hd, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h14, 8'h11, 8'hd, 8'h14, 8'h14, 8'hd, 8'hd, 8'h14, 8'h13, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h14, 8'h3, 8'hd, 8'h14, 8'h13, 8'h13, 8'h13, 8'h14, 8'h13, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h14, 8'h17, 8'hd, 8'h14, 8'h13, 8'h13, 8'h13, 8'h14, 8'h13, 8'h17, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h15, 8'h15, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h17, 8'h3, 8'h3, 8'h3, 8'h11, 8'he, 8'h15, 8'h15, 8'he, 8'he, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h6, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h3, 8'h12, 8'h15, 8'h15, 8'he, 8'h7, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h2, 8'h2, 8'h8, 8'h11, 8'h11, 8'h3, 8'h14, 8'h14, 8'h12, 8'h15, 8'h17, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'ha, 8'h2, 8'h11, 8'h11, 8'h3, 8'h13, 8'h13, 8'h17, 8'h17, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'ha, 8'h2, 8'h3, 8'h11, 8'h3, 8'hd, 8'h13, 8'hd, 8'h17, 8'h15, 8'h15, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h11, 8'h11, 8'h3, 8'h12, 8'h15, 8'h15, 8'hf, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h7, 8'h7, 8'h7, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};

ashRight0 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h7, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h11, 8'h15, 8'h15, 8'h1, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h7, 8'he, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h1, 8'h1, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'hd, 8'h13, 8'h13, 8'h3, 8'hd, 8'hd, 8'hd, 8'h11, 8'hd, 8'hd, 8'hd, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h14, 8'h14, 8'h17, 8'h13, 8'h13, 8'h13, 8'h11, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h14, 8'h14, 8'h13, 8'h13, 8'h14, 8'h14, 8'h3, 8'h14, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h14, 8'h14, 8'h13, 8'h13, 8'h14, 8'h14, 8'h17, 8'h14, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h17, 8'h17, 8'h1, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'hf, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h2, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'he, 8'hd, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h8, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h15, 8'he, 8'h17, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h2, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h15, 8'h15, 8'h11, 8'h11, 8'h3, 8'h13, 8'h13, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h11, 8'h11, 8'h3, 8'h13, 8'h13, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h17, 8'h17, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0 };
            ashRight1 = ' {8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'hf, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h15, 8'h3, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h15, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h15, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h1, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'hd, 8'h13, 8'h14, 8'h3, 8'hd, 8'h13, 8'hd, 8'hd, 8'h11, 8'h13, 8'h13, 8'h13, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h13, 8'h14, 8'hd, 8'h13, 8'h13, 8'h14, 8'h14, 8'h3, 8'h14, 8'hd, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'hf, 8'h13, 8'h13, 8'h14, 8'h13, 8'h13, 8'h13, 8'h14, 8'h12, 8'h17, 8'h14, 8'hd, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h17, 8'h11, 8'h15, 8'hd, 8'hd, 8'hd, 8'h13, 8'h13, 8'h13, 8'h14, 8'h13, 8'hd, 8'hd, 8'hd, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h11, 8'h15, 8'h17, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h15, 8'h15, 8'h15, 8'h17, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h15, 8'h15, 8'h15, 8'h17, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h17, 8'h15, 8'h15, 8'h15, 8'ha, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'hd, 8'h17, 8'h17, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h17, 8'he, 8'h7, 8'hd, 8'h8, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h14, 8'h14, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h3, 8'h11, 8'h11, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h13, 8'h13, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h15, 8'he, 8'h11, 8'h11, 8'h2, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'hd, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h15, 8'h7, 8'h11, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h3, 8'h1, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
ashRight2 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'hf, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h7, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h15, 8'h1, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h15, 8'h1, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h1, 8'h17, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h3, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h3, 8'h1, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h17, 8'h3, 8'h3, 8'h17, 8'h17, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h13, 8'h14, 8'h17, 8'h17, 8'h14, 8'h14, 8'h11, 8'h11, 8'h14, 8'h14, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h13, 8'h14, 8'h17, 8'h17, 8'h13, 8'h13, 8'h3, 8'h11, 8'h13, 8'h13, 8'hd, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h13, 8'h14, 8'h13, 8'h13, 8'h13, 8'h14, 8'h17, 8'h17, 8'h14, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h15, 8'he, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h7, 8'h15, 8'h15, 8'he, 8'h11, 8'h3, 8'h3, 8'h3, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h3, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'he, 8'he, 8'h15, 8'h15, 8'h12, 8'h3, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h15, 8'h12, 8'h14, 8'h14, 8'h11, 8'h11, 8'h11, 8'h2, 8'h2, 8'h2, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'he, 8'hd, 8'h14, 8'h14, 8'h11, 8'h11, 8'h11, 8'h2, 8'ha, 8'ha, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h15, 8'h15, 8'h17, 8'h1, 8'h13, 8'h13, 8'h11, 8'h11, 8'h11, 8'h8, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'hf, 8'he, 8'h15, 8'h12, 8'h3, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h7, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};

            ashUp0 = ' {8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h17, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h1, 8'h17, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h17, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h3, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h3, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h17, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h17, 8'h3, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h14, 8'h14, 8'h11, 8'h2, 8'h15, 8'h15, 8'h8, 8'h8, 8'h8, 8'h8, 8'h8, 8'h8, 8'h15, 8'h2, 8'ha, 8'h11, 8'h14, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h14, 8'h14, 8'h11, 8'h2, 8'h15, 8'h15, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h15, 8'h2, 8'ha, 8'h11, 8'h14, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h17, 8'h8, 8'h17, 8'h17, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h17, 8'h8, 8'ha, 8'h17, 8'h13, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h11, 8'h11, 8'he, 8'he, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'he, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h17, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h3, 8'h15, 8'h3, 8'h3, 8'h3, 8'h15, 8'h15, 8'h3, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
ashUp1 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h1, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h1, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h1, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h17, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h1, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h17, 8'h3, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h15, 8'h2, 8'h8, 8'h8, 8'h8, 8'h8, 8'h8, 8'h15, 8'h2, 8'h2, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'hd, 8'h17, 8'h11, 8'h2, 8'h2, 8'h17, 8'h5, 8'h5, 8'h5, 8'h5, 8'h5, 8'h5, 8'h17, 8'h2, 8'h2, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h13, 8'hd, 8'h11, 8'h2, 8'h2, 8'h17, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h3, 8'h2, 8'h2, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h13, 8'h13, 8'h13, 8'h8, 8'h2, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h2, 8'h8, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'hf, 8'h15, 8'h15, 8'hd, 8'hd, 8'h15, 8'h15, 8'hf, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h7, 8'h7, 8'h3, 8'h3, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h1, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
         ashUp2 = ' {8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h17, 8'h17, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h17, 8'h3, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h1, 8'h1, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h1, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h2, 8'h15, 8'hd, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'hd, 8'h15, 8'h3, 8'h3, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h2, 8'he, 8'hd, 8'h5, 8'h5, 8'h5, 8'h5, 8'h5, 8'hd, 8'h17, 8'h2, 8'h2, 8'h11, 8'h17, 8'hd, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h2, 8'h3, 8'h17, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h17, 8'h3, 8'h2, 8'h2, 8'h11, 8'h13, 8'h13, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h8, 8'he, 8'he, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'he, 8'he, 8'h8, 8'h8, 8'h17, 8'h13, 8'h13, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'ha, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'ha, 8'ha, 8'hd, 8'h1, 8'hd, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h15, 8'h15, 8'h15, 8'he, 8'h15, 8'he, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h3, 8'h3, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h7, 8'h15, 8'h17, 8'h17, 8'h17, 8'h15, 8'h7, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
end

logic [7:0] font_data;

logic [10:0] font_addr;
spriteROM sr0(.Sprite(pokemon_id), .frameClk(frameClk), .read_address(spriteAddr), .Clk(VGA_CLK), .data_Out(spriteData), .user_on(user_on), .pkmnID(userPokemonSprite), .wildPkmnID(wildPokemonSprite));

colorTable c0(.color(color), .DrawX(temp_X), .DrawY(temp_Y), .*);

font_rom f0(.addr(font_addr), .data(font_data));

logic wild1_on, wild2_on, wild3_on, wild4_on, wild5_on, wild6_on, wild7_on, wild8_on, wild9_on, wild10_on;
logic poke1_on, poke2_on, poke3_on, poke4_on, poke5_on, poke6_on, poke7_on, poke8_on, poke9_on, poke10_on;
logic level1_on, level2_on, level3_on, level4_on, level5_on, level6_on, level7_on, level8_on;
//Defining shape_on bits for font addressing for the pokemon names
always_comb
begin
//Setting default values
font_addr = 10'b0;
//pointer_on = 3'b000;
//
//poke_select1 = 1'b0;
//poke_select2 = 1'b0;
//poke_select3 = 1'b0;
            wild1_on = 1'b0;
wild2_on = 1'b0;
           wild3_on = 1'b0;
wild4_on = 1'b0;
           wild5_on = 1'b0;
wild6_on = 1'b0;
           wild7_on = 1'b0;
wild8_on = 1'b0;
           wild9_on = 1'b0;
wild10_on = 1'b0;
            poke1_on = 1'b0;
poke2_on = 1'b0;
           poke3_on = 1'b0;
poke4_on = 1'b0;
           poke5_on = 1'b0;
poke6_on = 1'b0;
           poke7_on = 1'b0;
poke8_on = 1'b0;
           poke9_on = 1'b0;
poke10_on = 1'b0;
            level1_on = 1'b0;
level2_on = 1'b0;
            level3_on = 1'b0;
level4_on = 1'b0;
            level5_on = 1'b0;
level6_on = 1'b0;
            level7_on = 1'b0;
level8_on = 1'b0;
            //Wild_pokemon Names
            if(DrawX >= 50 && DrawX < 58 && DrawY >= 25 && DrawY <=40)
            begin
            font_addr = (DrawY - 25 + 16*w[0]);//B
            wild1_on = 1'b1;
end


else if (DrawX >= 58 && DrawX < 66 && DrawY >= 25 && DrawY <= 40)
	begin
	font_addr = (DrawY - 25 + 16 * w[1]); //u
   wild2_on = 1'b1;
           end

           else if(DrawX >= 66 && DrawX < 74 && DrawY >= 25 && DrawY <=40)
           begin
           font_addr = (DrawY - 25 + 16*w[2]);//l
           wild3_on = 1'b1;
end


else if (DrawX >= 74 && DrawX < 82 && DrawY >= 25 && DrawY <= 40)
	begin
	font_addr = (DrawY - 25 + 16 * w[3]); //b
wild4_on = 1'b1;
           end

           else if(DrawX >= 82 && DrawX < 90 && DrawY >= 25 && DrawY <=40)
           begin
           font_addr = (DrawY - 25 + 16*w[4]);//a
           wild5_on = 1'b1;
end

else if (DrawX >= 90 && DrawX < 98 && DrawY >= 25 && DrawY <= 40)
	begin
	font_addr = (DrawY - 25 + 16 * w[5]); //s
wild6_on = 1'b1;
           end

           else if(DrawX >= 98 && DrawX < 106 && DrawY >= 25 && DrawY <=40)
           begin
           font_addr = (DrawY - 25 + 16*w[6]);//a
           wild7_on = 1'b1;
end

else if (DrawX >= 106 && DrawX < 114 && DrawY >= 25 && DrawY <= 40)
	begin
	font_addr = (DrawY - 25 + 16 * w[7]); //u
wild8_on = 1'b1;
           end


           else if(DrawX >= 114 && DrawX < 122 && DrawY >= 25 && DrawY <=40)
           begin
           font_addr = (DrawY - 25 + 16*w[8]);//r
           wild9_on = 1'b1;
end


else if (DrawX >= 122 && DrawX < 130 && DrawY >= 25 && DrawY <= 40)
	begin
	font_addr = (DrawY - 25 + 16 * w[9]); // WhiteSpace
wild10_on = 1'b1;
            end

            //User Pokemon Names
            else if(DrawX >= 310 && DrawX < 318 && DrawY >= 225 && DrawY <= 240)
            begin
            font_addr = (DrawY - 225 + 16*u[0]);//C
            poke1_on = 1'b1;
end

else if (DrawX >= 318 && DrawX < 326 && DrawY >= 225 && DrawY <= 240)
	begin
	font_addr = (DrawY - 225 + 16 * u[1]); //h
poke2_on = 1'b1;
           end

           else if(DrawX >= 326 && DrawX < 334 && DrawY >= 225 && DrawY <= 240)
           begin
           font_addr = (DrawY - 225 + 16*u[2]);//a
           poke3_on = 1'b1;
end

else if (DrawX >= 334 && DrawX < 342 && DrawY >= 225 && DrawY <= 240)
	begin
	font_addr = (DrawY - 225 + 16 * u[3]); //r
poke4_on = 1'b1;
           end

           else if(DrawX >= 342 && DrawX < 350 && DrawY >= 225 && DrawY <= 240)
           begin
           font_addr = (DrawY - 225 + 16*u[4]);//m
           poke5_on = 1'b1;
end

else if (DrawX >= 350 && DrawX < 358 && DrawY >= 225 && DrawY <= 240)
	begin
	font_addr = (DrawY - 225 + 16 * u[5]); //a
poke6_on = 1'b1;
           end

           else if(DrawX >= 358 && DrawX < 366 && DrawY >= 225 && DrawY <= 240)
           begin
           font_addr = (DrawY - 225 + 16*u[6]);//n
           poke7_on = 1'b1;
end

else if (DrawX >= 366 && DrawX < 374 && DrawY >= 225 && DrawY <= 240)
	begin
	font_addr = (DrawY - 225 + 16 * u[7]); //d
poke8_on = 1'b1;
           end

           else if(DrawX >= 374 && DrawX < 382 && DrawY >= 225 && DrawY <= 240)
           begin
           font_addr = (DrawY - 225 + 16*u[8]);//e
           poke9_on = 1'b1;
end


else if (DrawX >= 382 && DrawX < 390 && DrawY >= 225 && DrawY <= 240)
	begin
	font_addr = (DrawY - 225 + 16 * u[9]); //r
poke10_on = 1'b1;
            end

            else if(DrawX >= 560 && DrawX < 568 && DrawY >= 10 && DrawY <= 25)
            begin
            font_addr = (DrawY - 10 + 16*'h4c);//L
level1_on = 1'b1;
            end
            else if(DrawX >= 568 && DrawX < 576 && DrawY >= 10 && DrawY <= 25)
            begin
            font_addr = (DrawY - 10 + 16*'h65);//e
level2_on = 1'b1;
            end
            else if(DrawX >= 576 && DrawX < 584 && DrawY >= 10 && DrawY <= 25)
            begin
            font_addr = (DrawY - 10 + 16*'h76);//v
level3_on = 1'b1;
            end
            else if(DrawX >= 584 && DrawX < 592 && DrawY >= 10 && DrawY <= 25)
            begin
            font_addr = (DrawY - 10 + 16*'h65);//e
level4_on = 1'b1;
            end
            else if(DrawX >= 592 && DrawX < 600 && DrawY >= 10 && DrawY <= 25)
            begin
            font_addr = (DrawY - 10 + 16*'h6c);//l
level5_on = 1'b1;
            end
            else if(DrawX >= 600 && DrawX < 608 && DrawY >= 10 && DrawY <= 25)
            begin
            font_addr = (DrawY - 10 + 16*'h3a);//:
level6_on = 1'b1;
            end
            else if(DrawX >= 608 && DrawX < 616 && DrawY >= 10 && DrawY <= 25)
            begin
            font_addr = (DrawY - 10 + 16*'h00);//WhiteSpace --> Will be filled up
level7_on = 1'b1;
            end
            else if(DrawX >= 616 && DrawX < 624 && DrawY >= 10 && DrawY <= 25)
            begin
            font_addr = (DrawY - 10 + 16*'h35);//5
level8_on = 1'b1;
            end


            end

            //////////////////Uncomment from here//////////////////
            always_comb
            begin
				//pointer_on = 3'b100;
				//font_addr = 10'd0;
            curr_map = 2'b00;
				user_on = 1'b0;
color = 8'd35;
        pokemon_id = 2'b11; //This is set to 2'b11 so that no other pokemon sprites are loaded --> Make sure this is 2'b11 in all other stages except PokeSelect
spriteAddr = ((DrawY - 100) * 96) + (DrawX - ((pokemon_id + 1) * 150));
//display_control == 2'b00 --> INIT_STAGE
if (display_control == 2'b00)
        begin
        color = Data;
        end

        else if (display_control == 2'b01)  //POKE SELECT
begin
//pokemon_id = 2'b00;
//curr_map = 2'b01;
//pokemon_id = 2'b11;
//spriteAddr = ((DrawY-100)*96) + (DrawX - ((pokemon_id + 1)* 150));
//	if(keycode == 8'h04)
//   begin
//
//	end
//
//	else if(keycode == 8'h16)
//	begin
//
//	end
//
//	else if(keycode == 8'h07)
//	begin
//
//	end


if (DrawX >= 150 && DrawX < 246 && DrawY >= 100 && DrawY < 196)
	begin
	pokemon_id = 2'b00;
	             spriteAddr = ((DrawY-100)*96) + (DrawX - ((pokemon_id + 1)* 150));
	             if(spriteData == 8'h0)
	color = 8'd35;
	        else
	        color = spriteData;

	        end
	        else if(DrawX >= 300 && DrawX < 396 && DrawY >= 100 && DrawY < 196)
	        begin
	        pokemon_id = 2'b01;
	spriteAddr = ((DrawY - 100) * 96) + (DrawX - ((pokemon_id + 1) * 150));
	if (spriteData == 8'h0)
		        color = 8'd35;
		else
			color = spriteData;

			end
			else if (DrawX >= 450 && DrawX < 546 && DrawY >= 100 && DrawY < 196)
				begin
				pokemon_id = 2'b10;
				             spriteAddr = ((DrawY-100)*96) + (DrawX - ((pokemon_id + 1)* 150));
				             if(spriteData == 8'h0)
				color = 8'd35;
				        else
				        color = spriteData;

				        end
				        else
				        begin
				        //pokemon_id = 2'b11;
//spriteAddr = ((DrawY-100)*96) + (DrawX - ((pokemon_id + 1)* 150));
				color = 8'd35;

				        end



				        end

				        else if(display_control== 2'b10)  //MAP1 STAGE
				begin
				pokemon_id = 2'b11;
				             curr_map = 2'b01;
				spriteAddr = ((DrawY - 100) * 96) + (DrawX - ((pokemon_id + 1) * 150));
				if ( ( DistX >= 0 && DistX <= 28  && DistY >= 0 && DistY <= 40))


					begin

// Assign color based on ball_on signal



					if (ashDown0[DistY * 28 + DistX] != 8'h0 && spriteDirControl == 2'b00 && counter[3:2] == 2'b00  )
						        begin
						        color = ashDown0[DistY*28 +DistX];
						        end

						        else if (ashDown1[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b00 && counter[3:2] == 2'b01 )
						begin
						color = ashDown1[DistY * 28 + DistX];
						end

						else if (ashDown2[DistY * 28 + DistX] != 8'h0 && spriteDirControl == 2'b00 && counter[3:2] == 2'b10 )
							         begin
							         color = ashDown2[DistY*28 +DistX];
							         end

							         else if (ashLeft0[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b01 && counter[3:2] == 2'b00 )
							begin
							color = ashLeft0[DistY * 28 + DistX];
							end

							else if (ashLeft1[DistY * 28 + DistX] != 8'h0 && spriteDirControl == 2'b01 && counter[3:2] == 2'b01)
								         begin
								         color = ashLeft1[DistY*28 +DistX];
								         end

								         else if (ashLeft2[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b01 && counter[3:2] == 2'b10)
								begin
								color = ashLeft2[DistY * 28 + DistX];
								end

								else if (ashRight0[DistY * 28 + DistX] != 8'h0 && spriteDirControl == 2'b10 && counter[3:2] == 2'b00 )
									         begin
									         color = ashRight0[DistY*28 +DistX];
									         end

									         else if (ashRight1[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b10 && counter[3:2] == 2'b01)
									begin
									color = ashRight1[DistY * 28 + DistX];
									end

									else if (ashRight2[DistY * 28 + DistX] != 8'h0 && spriteDirControl == 2'b10 && counter[3:2] == 2'b10)
										         begin
										         color = ashRight2[DistY*28 +DistX];
										         end

										         else if (ashUp0[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b11 && counter[3:2] == 2'b00 )
										begin
										color = ashUp0[DistY * 28 + DistX];
										end

										else if (ashUp1[DistY * 28 + DistX] != 8'h0 && spriteDirControl == 2'b11 && counter[3:2] == 2'b01)
											         begin
											         color = ashUp1[DistY*28 +DistX];
											         end

											         else if (ashUp2[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b11 && counter[3:2] == 2'b10)
											begin
											color = ashUp2[DistY * 28 + DistX];
											end

											else if (ashDown0[DistY * 28 + DistX] == 8'h0|| ashDown1[DistY*28 +DistX]==8'h0 || ashDown2[DistY * 28 + DistX] == 8'h0|| ashLeft0[DistY*28 +DistX]==8'h0 || ashLeft1[DistY * 28 + DistX] == 8'h0|| ashLeft2[DistY*28 +DistX]==8'h0 || ashRight0[DistY * 28 + DistX] == 8'h0||ashRight1[DistY*28 +DistX]==8'h0 || ashRight2[DistY * 28 + DistX] == 8'h0|| ashUp0[DistY*28 +DistX]==8'h0 || ashUp1[DistY * 28 + DistX] == 8'h0||ashUp2[DistY*28 +DistX]==8'h0)

												begin

												color = Data;
												end

												end
												else
													begin
													if (level1_on == 1'b1 && font_data[560 - DrawX])
														        color = 8'd09;
														else if (level2_on == 1'b1 && font_data[568 - DrawX])
															         color = 8'd09;
															else if (level3_on == 1'b1 && font_data[576 - DrawX])
																         color = 8'd09;
																else if (level4_on == 1'b1 && font_data[584 - DrawX])
																	         color = 8'd09;
																	else if (level5_on == 1'b1 && font_data[592 - DrawX])
																		         color = 8'd09;
																		else if (level6_on == 1'b1 && font_data[600 - DrawX])
																			         color = 8'd09;
																			else if (level7_on == 1'b1 && font_data[608 - DrawX])
																				         color = 8'd09;
																				else if (level8_on == 1'b1 && font_data[616 - DrawX])
																					         color = 8'd09;
																					else
																						color = Data;
																						end



																						end


//////////////////Uncomment from here//////////////////
//
//		   else if( DrawX >= 42 && DrawX <= 146 && DrawY == 66 ) // Poke center top border
//		  begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawX >=42 && DrawX<=146 && DrawY== 146) //Poke center bottom border
//		  begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawY >=66 && DrawY<=146 && DrawX== 42) //Poke center left border
//		  begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawY >=66 && DrawY<=146 && DrawX== 146) //Poke center right border
//		  begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawX==0 && DrawY==30) // Left top corner of the map
//         begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawX==10 && DrawY==30) // Left top corner of the map
//         begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawX==20 && DrawY==30) // Left top corner of the map
//         begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawX==30 && DrawY==30) // Left top corner of the map
//         begin
//		  color = 8'd0;
//		  end
//
//		   else if(DrawX==0 && DrawY==480)    //Left bottom corner of the map
//         begin
//		  color = 8'd0;
//		  end
//
//		   else if(DrawX==640 && DrawY==0) // Right top corner
//         begin
//		  color = 8'd0;
//		  end

//		   else if(DrawX==640 && DrawY==480) // Right bottom
//         begin
//		  color = 8'd0;
//		  end




																						else if (display_control == 2'b11)
																							         begin
																							         pokemon_id = 2'b11;
																							curr_map = 2'b00;
																							           spriteAddr = ((DrawY - 50)*96 + (DrawX - 500));



																							           //Wild Pokemon Normal
																							           if(DrawX>= 500 && DrawX <= 596 && DrawY >= 50 && DrawY < 146 && battle_control != 4'b0110)
																							begin

																							spriteAddr = ((DrawY - 50) * 96 + (DrawX - 500));
																							if (spriteData == 8'h0)
																								        color = 8'd36;
																								else
																									color = spriteData;

																									end
//UserPokemon attacking
else if (DrawX >= 100 && DrawX < 196 && DrawY >= 250 && DrawY < 346 && battle_control == 4'b0011)
	   begin
spriteAddr = ((DrawY - 250)*96 + (DrawX - 100));
user_on = 1'b1;
 if(spriteData == 8'h0)
color = 8'd36;
else
color = spriteData;
end

//User Pokemon Normal
else if(DrawX >= 50 && DrawX <= 146 && DrawY >= 250 && DrawY < 346 && battle_control != 4'b0011)
begin
user_on = 1'b1;
spriteAddr = ((DrawY - 250) * 96 + DrawX - 50);
if (spriteData == 8'h0)
color = 8'd36;
else
color = spriteData;
end
else if (DrawX >= 450 && DrawX < 546 && DrawY >= 50 && DrawY < 146 && battle_control == 4'b0110)
begin
spriteAddr = ((DrawY - 50)*96 + (DrawX - 470));
if(spriteData == 8'h0)
color = 8'd36;
else
color = spriteData;
end
//Hp_WildPokemon Bar
else if(DrawX >= 50 && DrawX <= ((hp_poke2 * 4) + 50)  && DrawY >= 50 && DrawY <= 60)
begin
color = 8'd37;
spriteAddr =  ((DrawY - 250) * 96 + DrawX - 50);
end
//Hp_User_PokeBar
else if (DrawX >= 306 && DrawX <= ((hp_poke1 * 4) + 306)  && DrawY >= 250 && DrawY <= 260)
begin
color = 8'd37;
spriteAddr = ((DrawY - 250)*96 + DrawX - 50);
end
																															        //TextBox
else if((DrawX >= 0 && DrawX <= 639 && DrawY >= 340 && DrawY <= 345) || (DrawX >= 0 && DrawX <=5 && DrawY >= 340 && DrawY <= 479)|| (DrawX >= 629 && DrawX <=639 && DrawY >= 340 && DrawY <= 479)|| ((DrawX >= 0 && DrawX <=639 && DrawY >= 469 && DrawY <= 479)))
begin
color = 8'd09;
spriteAddr = ((DrawY - 250) * 96 + DrawX - 50);
end

else if (wild1_on == 1'b1 && font_data[58 - DrawX])
color = 8'd09;

else if (wild2_on == 1'b1 && font_data[66 - DrawX])
color = 8'd09;

else if (wild3_on == 1'b1 && font_data[74 - DrawX])
color = 8'd09;

else if (wild4_on == 1'b1 && font_data[82 - DrawX])
color = 8'd09;

else if (wild5_on == 1'b1 && font_data[90 - DrawX])
color = 8'd09;

else if (wild6_on == 1'b1 && font_data[98 - DrawX])
color = 8'd09;

else if (wild7_on == 1'b1 && font_data[106 - DrawX])
color = 8'd09;

else if (wild8_on == 1'b1 && font_data[114 - DrawX])
color = 8'd09;

else if (wild9_on == 1'b1 && font_data[122 - DrawX])
																																						                                                                    color = 8'd09;

																																						                                                                    else if (wild10_on == 1'b1 && font_data[130 - DrawX])
																																							                                                                            color = 8'd09;

																																							                                                                            else if (poke1_on == 1'b1 && font_data[318 - DrawX])
																																								                                                                                    color = 8'd09;

																																								                                                                                    else if (poke2_on == 1'b1 && font_data[326 - DrawX])
																																									                                                                                            color = 8'd09;

																																									                                                                                            else if (poke3_on == 1'b1 && font_data[334 - DrawX])
																																										                                                                                                    color = 8'd09;


																																										                                                                                                    else if (poke4_on == 1'b1 && font_data[342 - DrawX])
																																											                                                                                                            color = 8'd09;


																																											                                                                                                            else if (poke5_on == 1'b1 && font_data[350 - DrawX])
																																												                                                                                                                    color = 8'd09;


																																												                                                                                                                    else if (poke6_on == 1'b1 && font_data[358 - DrawX])
																																													                                                                                                                            color = 8'd09;


																																													                                                                                                                            else if (poke7_on == 1'b1 && font_data[366 - DrawX])
																																														                                                                                                                                    color = 8'd09;


																																														                                                                                                                                    else if (poke8_on == 1'b1 && font_data[374 - DrawX])
																																															                                                                                                                                            color = 8'd09;


																																															                                                                                                                                            else if (poke9_on == 1'b1 && font_data[382 - DrawX])
																																																                                                                                                                                                    color = 8'd09;


																																																                                                                                                                                                    else if (poke10_on == 1'b1 && font_data[390 - DrawX])
																																																	                                                                                                                                                            color = 8'd09;






//Background for battle --> Make it load from SRAM
else
begin
color = 8'd36;
spriteAddr = ((DrawY - 250)*96 + DrawX - 50);
end

end

end
endmodule




																																																		                                                                                                                                                                    // NOTE: add curr_map_pixel



																																																		                                                                                                                                                                    //logic ball_on;


																																																		                                                                                                                                                                    //
																																																		                                                                                                                                                                    //logic ash_on;
																																																		                                                                                                                                                                    //logic [7:0] Red, Green, Blue;
																																																		                                                                                                                                                                    //
																																																		                                                                                                                                                                    //
																																																		                                                                                                                                                                    //
																																																		                                                                                                                                                                    ///* The ball's (pixelated) circle is generated using the standard circle formula.  Note that while
//   the single line is quite powerful descriptively, it causes the synthesis tool to use up three
//   of the 12 available multipliers on the chip! Since the multiplicants are required to be signed,
//   we have to first cast them from logic to int (signed by default) before they are multiplied. */
//
//int DistX, DistY, Size;
//assign DistX = DrawX - BallX;
//assign DistY = DrawY - BallY;
////assign Size = BallS;
//
//assign VGA_R = Red;
//assign VGA_G = Green;
//assign VGA_B = Blue;
//
////logic [7:0] MAP1[0:76799];
////logic [15:0] curr_map_pixel;
//
//
//logic [7:0] ashDown0[0:1119];
//logic [7:0] ashDown1[0:1119];
//logic [7:0] ashDown2[0:1119];
//
//logic [7:0] ashLeft0[0:1119];
//logic [7:0] ashLeft1[0:1119];
//logic [7:0] ashLeft2[0:1119];
//
//logic [7:0] ashRight0[0:1119];
//logic [7:0] ashRight1[0:1119];
//logic [7:0] ashRight2[0:1119];
//
//logic [7:0] ashUp0[0:1119];
//logic [7:0] ashUp1[0:1119];
//logic [7:0] ashUp2[0:1119];
//
//
//logic [15:0] color;
//logic [1:0] pokemon_id;
//logic [7:0] spriteData;
//logic [13:0] spriteAddr;
//
//
////logic [10:0] font_addr;
////logic [7:0] font_data;
////
////logic [9:0] temp_X, temp_Y;
////assign temp_X = DrawX;
////assign temp_Y = DrawY;
//
////logic [7:0] temp;
//
//always_comb
//begin
//
//if(DrawX >= 150 && DrawX <216 && DrawY >= 100 && DrawY < 196)
//begin
//pokemon_id = 2'b00;
//
//end
//else if(DrawX >= 300 && DrawX < 396 && DrawY >= 100 && DrawY < 196)
//begin
//pokemon_id = 2'b01;
////spriteAddr = (DrawY-100) * 96 + (DrawX - 240);
//end
//else if(DrawX >= 450 && DrawX < 546 && DrawY >= 100 && DrawY < 196)
//begin
//pokemon_id = 2'b10;
////spriteAddr = (DrawY-100) * 96 + (DrawX - 360);
//end
//else
//pokemon_id = 2'b11;
////spriteAddr = 0;
//end
////assign pixel = (DrawY/2) * 320 + (DrawX/2);
//assign spriteAddr = ((DrawY-100)*96) + (DrawX - ((pokemon_id + 1)* 150));
//
//spriteROM sr0(.Sprite(pokemon_id), .read_address(spriteAddr), .Clk(Clk), .data_Out(spriteData));
//
//always_comb
//begin
//
//if((pokemon_id == 2'b00 || pokemon_id == 2'b01 || pokemon_id == 2'b10) && spriteData != 8'h0)
//begin
//temp = 0;
//color = spriteData;
////font_addr = 16*'h0;
//end
//else if(DrawX >= 150 && DrawX <= 450 && DrawY >= 400 && DrawY <= 420)
//begin
//temp = 0;
//if(DrawX>= 150 && DrawX <= 160 && DrawY >= 400 && DrawY <= 420)
//begin
//temp = 16*'h50;
//if(font_addr[DrawX - 150] == 1'b1)
//color = 8'd17;
//else
//color = 8'd34;
//end
//else
//color = 8'd34;
//end
//
//
//
//
//else
//begin
////font_addr = 16*'h0;
//temp = 0;
//color = 8'd34;
//end
//end
//assign font_addr = 16*temp;
//
//font_rom font(.addr(font_addr), .data(font_data));
//
//colorTable c0(.color(color), .DrawX(temp_X), .DrawY(temp_Y), .*);

																																																			                                                                                                                                                                    /*
																																																			                                                                                                                                                                    always_ff
																																																			                                                                                                                                                                    					begin

																																																			                                                                                                                                                                              //MAP1 = '{ 8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'hd,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h16,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h16,8'hd,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'h1,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h1,8'h1,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h1,8'hb,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'h1,8'hd,8'h4,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h14,8'hc,8'h1,8'hd,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'h14,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'h14,8'h14,8'hc,8'h1,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'h14,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h6,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'h1,8'h14,8'h14,8'hc,8'h1,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'h14,8'h13,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'ha,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h14,8'h14,8'hc,8'h1,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'hb,8'h13,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'h13,8'h14,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'hd,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'h13,8'hd,8'hd,8'hd,8'hd,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hd,8'hd,8'h13,8'h1,8'hd,8'h17,8'ha,8'ha,8'h17,8'h17,8'ha,8'ha,8'h17,8'h17,8'hd,8'h13,8'hd,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'hb,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hd,8'h1,8'h17,8'h17,8'ha,8'ha,8'h17,8'h17,8'hd,8'hd,8'h17,8'h17,8'h17,8'ha,8'h17,8'h17,8'h17,8'hd,8'hd,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'hb,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'h1,8'h17,8'ha,8'h17,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'h17,8'ha,8'h17,8'h16,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'hb,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'h16,8'ha,8'ha,8'h17,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h1,8'h17,8'ha,8'h1,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'hc,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h14,8'hc,8'h1,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h13,8'h13,8'hb,8'h1,8'h17,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h1,8'h17,8'h1,8'hb,8'h13,8'h13,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'h1,8'hd,8'h9,8'hb,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h14,8'h14,8'h13,8'h1,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h16,8'h1,8'h4,8'h13,8'h14,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h14,8'h4,8'h13,8'h1,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h14,8'hc,8'hc,8'h4,8'h13,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h16,8'h1,8'h4,8'h14,8'h14,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h10,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h13,8'h4,8'h13,8'hc,8'h13,8'h16,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hc,8'h9,8'h9,8'h9,8'h9,8'h9,8'h13,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h16,8'h4,8'h4,8'h14,8'h4,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h1,8'h4,8'h4,8'h13,8'h14,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hc,8'h9,8'h4,8'h4,8'h13,8'h4,8'h9,8'h9,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'hb,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h14,8'h14,8'h14,8'hc,8'h13,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h1,8'hd,8'h4,8'h4,8'h14,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h4,8'h4,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h14,8'h13,8'hc,8'hc,8'h13,8'h13,8'h14,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h4,8'h4,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h14,8'hc,8'h13,8'h1,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h1,8'h1,8'h1,8'h4,8'h4,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h14,8'hc,8'h9,8'h9,8'h4,8'h13,8'h13,8'h13,8'h13,8'h13,8'h1,8'h1,8'h13,8'h9,8'h9,8'h4,8'h1,8'h1,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h9,8'h9,8'h9,8'h14,8'h13,8'hb,8'hb,8'hb,8'hb,8'h13,8'hc,8'h13,8'h1,8'h1,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h1,8'h1,8'h1,8'hd,8'h14,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'hc,8'h9,8'hc,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h4,8'h4,8'h13,8'h4,8'h4,8'h13,8'h4,8'h4,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h4,8'h9,8'h9,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h13,8'h1,8'h1,8'h1,8'h1,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h1,8'h1,8'h1,8'h1,8'hd,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h4,8'h9,8'h9,8'h4,8'h4,8'hc,8'h9,8'hc,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h1,8'h1,8'h1,8'h1,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h4,8'h9,8'h9,8'h9,8'h9,8'h4,8'hd,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'hd,8'h4,8'h4,8'hd,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h17,8'hd,8'hd,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hd,8'hd,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'hd,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'hd,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h1,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'hd,8'h10,8'ha,8'hd,8'h10,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'h4,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hd,8'h5,8'hd,8'h16,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hd,8'h5,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hc,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hc,8'hc,8'h4,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h1,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h16,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h4,8'hc,8'h9,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h10,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hc,8'hc,8'hc,8'h4,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h1,8'h16,8'h16,8'h16,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h16,8'h16,8'h16,8'h1,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hc,8'hc,8'h9,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hc,8'hc,8'hc,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'hd,8'ha,8'ha,8'hd,8'ha,8'h17,8'h17,8'h17,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h17,8'h17,8'h17,8'h17,8'hd,8'ha,8'ha,8'hd,8'h5,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'hc,8'hc,8'h9,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'h4,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hd,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'hc,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'ha,8'h4,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hd,8'ha,8'ha,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h4,8'hd,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'ha,8'ha,8'h4,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hd,8'ha,8'ha,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h10,8'ha,8'ha,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'hd,8'ha,8'ha,8'h4,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hd,8'ha,8'ha,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h5,8'ha,8'hd,8'hd,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'ha,8'hd,8'ha,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'hd,8'ha,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'ha,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'ha,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h4,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'ha,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'h7,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'h7,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'ha,8'ha,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h5,8'h5,8'h5,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'h5,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h7,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'h7,8'h5,8'h5,8'h5,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h5,8'h5,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'h5,8'h7,8'ha,8'ha,8'h11,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'ha,8'hf,8'ha,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h7,8'h5,8'hf,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'ha,8'h7,8'hf,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'ha,8'h11,8'ha,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h5,8'hf,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h7,8'h5,8'h7,8'hf,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'ha,8'ha,8'h11,8'h5,8'ha,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'h7,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'hf,8'ha,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'ha,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h11,8'ha,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'ha,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'h17,8'hd,8'h4,8'h10,8'h5,8'h10,8'h5,8'h4,8'hd,8'h17,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'h7,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'h7,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'h7,8'hf,8'h11,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'h17,8'h17,8'h17,8'hd,8'h4,8'h7,8'h7,8'h7,8'h7,8'h5,8'hd,8'h17,8'h17,8'h17,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h11,8'ha,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'ha,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'h17,8'h17,8'h17,8'h17,8'h17,8'hd,8'h4,8'hd,8'h7,8'h7,8'h7,8'h10,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'h17,8'h17,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'hd,8'h1,8'hd,8'hd,8'hd,8'hd,8'h17,8'h17,8'h7,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'h11,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'ha,8'h7,8'h7,8'h17,8'h17,8'h17,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'h17,8'h17,8'h7,8'h7,8'h7,8'ha,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h10,8'h10,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'ha,8'h7,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h7,8'ha,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'ha,8'h10,8'h5,8'h5,8'h5,8'h10,8'ha,8'h7,8'h11,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'h7,8'hd,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h13,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h10,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h10,8'h10,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h10,8'h10,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h3,8'h5,8'h10,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h10,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h17,8'hd,8'hd,8'hd,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h1,8'h1,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h7,8'ha,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'ha,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'ha,8'hf,8'hf,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h10,8'h5,8'ha,8'h5,8'h7,8'hf,8'ha,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'h7,8'h7,8'hf,8'h7,8'h3,8'h5,8'h5,8'h5,8'h10,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h3,8'h17,8'h17,8'h17,8'h17,8'h3,8'ha,8'h11,8'ha,8'ha,8'h11,8'ha,8'ha,8'h11,8'ha,8'h3,8'h1,8'hd,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h17,8'h17,8'h17,8'h17,8'h1,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h1,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h17,8'h3,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h3,8'h17,8'h17,8'hd,8'h5,8'hd,8'h5,8'h5,8'hd,8'h5,8'hd,8'hd,8'h5,8'hd,8'h17,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h1,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'hd,8'hd,8'hd,8'hd,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'hd,8'h1,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h17,8'h7,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'hd,8'hd,8'hd,8'h5,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h10,8'hd,8'h17,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h17,8'h7,8'ha,8'he,8'he,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h17,8'h17,8'hd,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hd,8'h17,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'h7,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h1,8'h7,8'ha,8'h17,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'hd,8'hd,8'hd,8'h4,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h4,8'hd,8'hd,8'h17,8'hd,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h11,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'h11,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h1,8'hd,8'h17,8'h17,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h1,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h17,8'h17,8'h17,8'h1,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h17,8'h17,8'h17,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'h17,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h7,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h7,8'h7,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'ha,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h7,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'h7,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h10,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h10,8'h5,8'h7,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h10,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'h7,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h10,8'h5,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'h7,8'hf,8'h11,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h11,8'ha,8'h10,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h7,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'h7,8'hf,8'h11,8'h7,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'ha,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h11,8'h11,8'ha,8'h7,8'ha,8'h10,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'h7,8'hf,8'ha,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h11,8'ha,8'h7,8'h7,8'h10,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'h11,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'ha,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'h11,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'ha,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'ha,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'ha,8'hf,8'hf,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hc,8'hc,8'h5,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h10,8'hc,8'hc,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h7,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h5,8'h8,8'hc,8'hc,8'h10,8'hd,8'ha,8'ha,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'ha,8'h5,8'hc,8'hc,8'h10,8'h8,8'hd,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h5,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h5,8'h7,8'hf,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h5,8'h5,8'hf,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'h5,8'hf,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h5,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h5,8'ha,8'hf,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'ha,8'h5,8'hf,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h5,8'hf,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h4,8'h4,8'hc,8'h10,8'hc,8'h10,8'ha,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'ha,8'ha,8'hc,8'hc,8'h10,8'h4,8'h4,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h7,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h7,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'h14,8'h4,8'h10,8'hc,8'h5,8'ha,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'h10,8'hc,8'h10,8'h4,8'h4,8'h10,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h4,8'h4,8'hc,8'h10,8'hc,8'h5,8'ha,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'hc,8'hc,8'h10,8'hc,8'h14,8'h4,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h12,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h14,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h14,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h14,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'ha,8'hf,8'h11,8'h7,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'h7,8'h7,8'h11,8'h7,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'ha,8'hf,8'h7,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'ha,8'hf,8'hf,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'h7,8'h7,8'h11,8'h7,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'h11,8'h7,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'ha,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h11,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h14,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'h7,8'h7,8'h10,8'h10,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'ha,8'h10,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h10,8'h10,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'h7,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h12,8'h4,8'h10,8'h10,8'hc,8'h5,8'ha,8'ha,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'ha,8'h10,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h10,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h10,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h14,8'h4,8'h10,8'h10,8'hc,8'h10,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hc,8'hc,8'h8,8'hc,8'h14,8'h4,8'h5,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h10,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'ha,8'h10,8'h10,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h10,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'hc,8'hc,8'h10,8'h8,8'h10,8'hc,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h4,8'h4,8'h4,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'hc,8'hc,8'h8,8'h8,8'hc,8'hc,8'hc,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hc,8'h4,8'h4,8'hc,8'h10,8'h8,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h9,8'h9,8'h9,8'h9,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h8,8'h8,8'hc,8'hc,8'h4,8'hc,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'h11,
																																																			                                                                                                                                                                              //8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h4,8'h4,8'h4,8'hc,8'h10,8'h8,8'h8,8'h8,8'h8,8'h10,8'h9,8'h9,8'hc,8'hc,8'hc,8'h9,8'h9,8'h10,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'hc,8'h9,8'h4,8'h4,8'h4,8'h2,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h2,8'h5,8'hc,8'h4,8'h12,8'hc,8'hc,8'hc,8'hc,8'h10,8'h10,8'hc,8'h10,8'h10,8'hc,8'hc,8'h10,8'hc,8'h10,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'hc,8'hc,8'hc,8'hc,8'h4,8'h12,8'hc,8'hc,8'h8,8'h2,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'h11,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'h11,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'hf,8'ha,8'h11,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'h11,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h2,8'h8,8'hc,8'h4,8'h14,8'h14,8'h4,8'h9,8'h10,8'h2,8'h2,8'h2,8'hc,8'h9,8'hc,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h4,8'h9,8'h9,8'h4,8'h14,8'h12,8'hc,8'hc,8'h8,8'h2,8'h2,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'h7,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'ha,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h2,8'h8,8'h2,8'h8,8'h8,8'hc,8'h4,8'h4,8'h9,8'h9,8'h10,8'h5,8'hc,8'h10,8'h10,8'h9,8'h4,8'h10,8'hc,8'h10,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'hc,8'h9,8'hc,8'h4,8'h4,8'hc,8'h8,8'h8,8'h2,8'h8,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h2,8'h8,8'h2,8'h8,8'h5,8'h10,8'h10,8'h10,8'h10,8'h5,8'h10,8'h9,8'h9,8'hc,8'h10,8'hc,8'h9,8'h9,8'h4,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'h10,8'h10,8'h10,8'h10,8'h8,8'h8,8'h2,8'h8,8'h2,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'hc,8'h9,8'h9,8'h9,8'h9,8'h9,8'hc,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'hd,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'ha,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'h5,8'h2,8'h8,8'h2,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h10,8'hc,8'hc,8'hc,8'h10,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h5,8'hd,8'hd,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'hd,8'h17,8'h5,8'h5,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h13,8'h17,8'h5,8'h5,8'hd,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hd,8'h5,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h5,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h2,8'h5,8'h5,8'hd,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h5,8'h7,8'hf,8'h7,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'h7,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'h5,8'hf,8'hf,8'h7,8'hf,8'h11,8'h11,8'h3,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'h7,8'hf,8'h7,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'ha,8'ha,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'hf,8'hf,8'h7,8'hf,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'h7,8'hf,8'h7,8'hf,8'h11,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h13,8'hd,8'h17,8'hd,8'hd,8'hd,8'hd,8'h10,8'h5,8'h5,8'h5,8'hd,8'h12,8'h12,8'hd,8'h17,8'h17,8'hd,8'h13,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'hd,8'hd,8'h17,8'hd,8'h13,8'hd,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'ha,8'hd,8'h5,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'h10,8'hd,8'hd,8'hd,8'hd,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h10,8'h10,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'ha,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h11,8'h7,8'h7,8'ha,8'h10,8'h5,8'h5,8'h10,8'h5,8'ha,8'h5,8'h7,8'h7,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'h5,8'ha,8'h7,8'h7,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h11,8'h7,8'h7,8'h7,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'h17,8'h4,8'h4,8'h4,8'h17,8'h5,8'h10,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'h17,8'hd,8'h4,8'h4,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h17,8'h17,8'h17,8'hd,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'h5,8'ha,8'hd,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'ha,8'hc,8'h4,8'ha,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h5,8'h10,8'h5,8'h5,8'ha,8'hf,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h10,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h10,8'h10,8'h5,8'ha,8'ha,8'hf,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'hd,8'h12,8'h13,8'hd,8'h17,8'ha,8'h10,8'h10,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h13,8'h12,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h4,8'h13,8'hd,8'h17,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'hc,8'h4,8'hd,8'h2,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h2,8'hd,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hc,8'h9,8'h4,8'ha,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'h7,8'h7,8'h7,8'h5,8'h10,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'h11,8'hf,8'hf,8'ha,8'h7,8'h5,8'h5,8'h5,8'h7,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h10,8'ha,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'ha,8'ha,8'h5,8'h7,8'hf,8'hf,8'h11,8'hf,8'ha,8'h7,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h13,8'hd,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'h17,8'h13,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'hc,8'hc,8'h4,8'ha,8'h5,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hc,8'h9,8'h9,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'h4,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'h4,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hc,8'hc,8'hc,8'h4,8'ha,8'h2,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h2,8'ha,8'ha,8'ha,8'ha,8'hd,8'h10,8'h10,8'h10,8'h10,8'h10,8'h5,8'h4,8'hc,8'hc,8'h9,8'h4,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'h11,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h3,8'hd,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h17,8'h13,8'h4,8'hd,8'h17,8'h3,8'h17,8'h4,8'hd,8'h17,8'hd,8'h5,8'h5,8'hd,8'hd,8'h4,8'h13,8'h17,8'h17,8'h17,8'h4,8'h4,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hc,8'hc,8'hc,8'hd,8'ha,8'ha,8'hd,8'ha,8'ha,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'ha,8'ha,8'hd,8'h2,8'ha,8'hd,8'ha,8'ha,8'hd,8'h10,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h5,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h17,8'h17,8'h4,8'h4,8'hd,8'h3,8'ha,8'h5,8'h5,8'hd,8'h17,8'hd,8'h17,8'h17,8'h3,8'hd,8'h4,8'hd,8'h17,8'h17,8'h5,8'h5,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'hd,8'h4,8'h13,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'h4,8'hc,8'hc,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h5,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h5,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'h11,8'h7,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'h11,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'h7,8'h11,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'hf,8'hf,8'h11,8'h7,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'ha,8'hf,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h17,8'hd,8'hd,8'h17,8'hd,8'hd,8'h17,8'h3,8'hd,8'h5,8'h5,8'h5,8'h17,8'h3,8'hd,8'hd,8'h17,8'hd,8'hd,8'h17,8'h3,8'h17,8'h5,8'h5,8'h5,8'ha,8'h3,8'h17,8'h13,8'h17,8'hd,8'hd,8'h17,8'h3,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'ha,8'h4,8'hc,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h5,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h9,8'h5,8'ha,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h11,8'hf,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h11,8'h11,8'h7,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'h7,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'hf,8'hf,8'h7,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h17,8'ha,8'hd,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h17,8'ha,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'ha,8'ha,8'hd,8'h17,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'ha,8'ha,8'h4,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h5,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'h5,8'ha,8'ha,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'h7,8'hf,8'hf,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'ha,8'hd,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'hd,8'h5,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hd,8'ha,8'hd,8'hd,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'h11,8'hf,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'ha,8'hd,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'hd,8'ha,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h11,8'h11,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hf,8'hf,8'h11,8'h11,8'h11,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'hd,8'ha,8'ha,8'ha,8'ha,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'ha,8'ha,8'ha,8'ha,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h13,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h13,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h13,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'hc,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'ha,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'ha,8'hf,8'h7,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'ha,8'h5,8'h5,8'h5,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'hf,8'h11,8'h7,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h5,8'h5,8'h5,8'h5,8'hf,8'h7,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'h12,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'hd,8'h17,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h10,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'h13,8'hd,8'h17,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'hd,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'h7,8'h5,8'ha,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'ha,8'h5,8'h5,8'h7,8'h5,8'h5,8'ha,8'h5,8'ha,8'hf,8'hf,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'hf,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h5,8'h5,8'ha,8'h5,8'h7,8'hf,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h17,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h17,8'h13,8'h4,8'h13,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'h17,8'h5,8'h5,8'h5,8'h10,8'h5,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h10,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'hc,8'h9,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'h6,8'h7,8'h10,8'h5,8'h5,8'h5,8'ha,8'ha,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h10,8'ha,8'h7,8'h7,8'h5,8'h10,8'h10,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h10,8'ha,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h17,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h10,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h10,8'h10,8'h5,8'h5,8'hd,8'hd,8'h17,8'h17,8'h13,8'h4,8'h12,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h10,8'h5,8'h17,8'hd,8'h17,8'h17,8'h4,8'h4,8'h13,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h17,8'hd,8'h17,8'h17,8'h4,8'h4,8'hd,8'h17,8'h5,8'h5,8'h10,8'h5,8'h5,8'hd,8'hd,8'h17,8'h17,8'h13,8'h4,8'h12,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'hd,8'h4,8'h4,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h6,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'ha,8'h7,8'h6,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h7,8'h6,8'h6,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'hd,8'hd,8'hd,8'h17,8'h13,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h13,8'hd,8'h17,8'h3,8'h5,8'h10,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'hd,8'h13,8'hd,8'hd,8'h17,8'ha,8'h10,8'h10,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'h13,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'h13,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'h13,8'hd,8'h17,8'h3,8'h5,8'h5,8'h10,8'h10,8'hd,8'hd,8'hd,8'hd,8'hd,8'h13,8'hd,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'hd,8'h13,8'hd,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'hd,8'h13,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'hd,8'h17,8'hd,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h4,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h6,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'ha,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h10,8'h5,8'h5,8'h10,8'h5,8'ha,8'h5,8'ha,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'h12,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h5,8'h10,8'h5,8'hd,8'h4,8'h4,8'h4,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'hd,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'h4,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'h4,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'hd,8'h13,8'h4,8'h4,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'hd,8'h5,8'h5,8'hd,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h5,8'ha,8'h7,8'h6,8'h6,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'ha,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h13,8'h4,8'h4,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'ha,8'h5,8'h5,8'hd,8'hd,8'h4,8'h4,8'hd,8'h17,8'h3,8'hd,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h3,8'hd,8'h12,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'h4,8'h17,8'h3,8'h17,8'h13,8'hd,8'h17,8'hd,8'h5,8'h5,8'hd,8'h13,8'h4,8'h4,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h3,8'hd,8'h13,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h4,8'h4,8'h13,8'h17,8'h3,8'h17,8'h12,8'hd,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'hd,8'h4,8'h4,8'hd,8'h17,8'h3,8'hd,8'h12,8'hd,8'h17,8'h5,8'h5,8'h5,8'h17,8'h4,8'h4,8'h4,8'h17,8'h17,8'h17,8'hd,8'hd,8'h17,8'hd,8'h5,8'h5,8'hd,8'hd,8'h4,8'h4,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'hd,8'h13,8'hd,8'h17,8'h3,8'hd,8'h4,8'h4,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h13,8'hd,8'h17,8'h17,8'h17,8'h4,8'h4,8'h17,8'h3,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h17,8'h17,8'h4,8'h4,8'hd,8'h3,8'hd,8'h5,8'h5,8'h17,8'hd,8'h13,8'h17,8'h17,8'h3,8'hd,8'h4,8'h13,8'h17,8'ha,8'h5,8'h5,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'hd,8'h4,8'h4,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h17,8'h17,8'h4,8'h4,8'hd,8'h3,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h17,8'h3,8'h4,8'h4,8'hd,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h17,8'h17,8'h4,8'h4,8'hd,8'h3,8'hd,8'h5,8'h5,8'h17,8'hd,8'h13,8'h17,8'h17,8'h3,8'hd,8'h4,8'h13,8'h17,8'h17,8'h5,8'h5,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'hd,8'h4,8'h4,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'h13,8'h17,8'hd,8'h13,8'hd,8'h3,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'hd,8'h17,8'hd,8'h12,8'hd,8'h17,8'h3,8'h5,8'h5,8'h5,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'hd,8'h17,8'hd,8'h13,8'h17,8'h3,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'h13,8'h17,8'hd,8'h13,8'hd,8'h3,8'h17,8'h5,8'h5,8'h5,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'h5,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hd,8'h17,8'h17,8'hd,8'hd,8'h17,8'h13,8'hd,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'hd,8'h17,8'hd,8'h13,8'h17,8'h3,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h17,8'h13,8'h17,8'hd,8'h13,8'hd,8'h3,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'hd,8'hd,8'h17,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'h17,8'h5,8'h5,8'h5,8'h5,8'h5,8'h17,8'hd,8'h17,8'h17,8'h17,8'h17,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'ha,8'hd,8'hd,8'h17,8'h17,8'hd,8'h17,8'h17,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'hd,8'h17,8'hd,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h7,8'h17,8'h7,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'hd,8'h17,8'h7,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'h7,8'h17,8'h7,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'h7,8'h17,8'h7,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h7,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'hd,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h17,8'h17,8'hd,8'h5,8'h5,8'h7,8'h17,8'h7,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h7,8'h17,8'hd,8'h5,8'h5,8'hd,8'h17,8'h7,8'h5,8'h5,8'h5,8'h17,8'h17,8'h5,8'h5,8'h5,8'h7,8'h17,8'h5,8'h5,8'h5,8'hd,8'h17,8'hd,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'h7,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'h7,8'h17,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'h5,8'h17,8'hd,8'h17,8'ha,8'h5,8'h17,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h17,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'ha,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'ha,8'h5,8'hd,8'h13,8'h13,8'h7,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'ha,8'h5,8'hd,8'h12,8'hd,8'h7,8'h5,8'h17,8'h13,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'h5,8'ha,8'hd,8'h12,8'hd,8'h7,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'hd,8'h5,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'ha,8'h5,8'hd,8'h13,8'hd,8'h7,8'h5,8'h17,8'h13,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'h5,8'h5,8'hd,8'h12,8'hd,8'h7,8'h5,8'h17,8'h13,8'h12,8'h17,8'h5,8'h7,8'hd,8'h12,8'hd,8'h5,8'ha,8'hd,8'h12,8'hd,8'h7,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'hd,8'h5,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h17,8'h13,8'h13,8'h17,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h17,8'h5,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h3,8'h5,8'h5,8'h17,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'hd,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h17,8'h5,8'h5,8'h3,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'h7,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'h7,8'h17,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h3,8'hd,8'hd,8'h7,8'h5,8'h7,8'hd,8'hd,8'h3,8'h5,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h10,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h17,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h17,8'h5,8'h17,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h17,8'h5,8'h17,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h17,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h17,8'h5,8'h17,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'h5,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h7,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h3,8'h3,8'h3,8'h3,8'hd,8'h17,8'h3,8'h3,8'h3,8'h7,8'ha,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'ha,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'h7,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'ha,8'ha,8'h3,8'h3,8'h3,8'h7,8'ha,8'h3,8'h3,8'h3,8'h3,8'hd,8'h3,8'h3,8'h3,8'h3,8'hd,8'h17,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h3,8'h3,8'h3,8'h3,8'hd,8'h7,8'h3,8'h3,8'h3,8'ha,8'ha,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h7,8'h3,8'h3,8'h3,8'hd,8'hd,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h17,8'h3,8'h3,8'h3,8'hd,8'hd,8'h3,8'h3,8'h3,8'h7,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h3,8'h3,8'h3,8'h3,8'hd,8'h7,8'h3,8'h3,8'h3,8'h7,8'hd,8'h3,8'h3,8'h3,8'h3,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'ha,8'h5,8'h7,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h3,8'ha,8'ha,8'ha,8'ha,8'h17,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h7,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h17,8'h7,8'h17,8'h17,8'h17,8'h5,8'h5,8'hd,8'h17,8'h17,8'h17,8'hd,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'ha,8'hd,8'h12,8'hd,8'ha,8'h5,8'h5,8'h17,8'hd,8'h13,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h10,8'hc,8'h9,8'h10,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'ha,8'hd,8'h13,8'hd,8'ha,8'h5,8'h5,8'h17,8'hd,8'h13,8'h17,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'ha,8'h3,8'hd,8'h3,8'ha,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'h5,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'ha,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'ha,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h5,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h10,8'ha,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'ha,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'ha,8'h3,8'hd,8'h3,8'ha,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'h5,8'ha,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'hd,8'h12,8'hd,8'h7,8'h5,8'h5,8'h17,8'hd,8'h12,8'h17,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'h17,8'h13,8'h17,8'h7,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'ha,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'ha,8'h3,8'h17,8'h3,8'h7,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h17,8'h13,8'h17,8'ha,8'h10,8'h5,8'h3,8'hd,8'hd,8'h3,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'ha,8'hd,8'h13,8'hd,8'h7,8'h5,8'h5,8'h17,8'hd,8'h12,8'h17,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'ha,8'h17,8'hd,8'h17,8'h3,8'h5,8'h5,8'h3,8'hd,8'hd,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'ha,8'h3,8'h3,8'h3,8'h7,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'ha,8'h17,8'h17,8'h17,8'ha,8'h10,8'h5,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'ha,8'hd,8'h13,8'hd,8'ha,8'h5,8'h5,8'h17,8'hd,8'h12,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'ha,8'h17,8'hd,8'h17,8'h7,8'h5,8'h5,8'h3,8'hd,8'hd,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'hc,8'h9,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'h3,8'h3,8'h3,8'h7,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'hc,8'h9,8'h5,8'h5,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'ha,8'h17,8'hd,8'h17,8'ha,8'h5,8'h5,8'h3,8'hd,8'hd,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'hd,8'h12,8'hd,8'h7,8'h5,8'h5,8'h3,8'hd,8'h13,8'h17,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h10,8'hc,8'h9,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'ha,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'hd,8'h3,8'h7,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h10,8'hc,8'h9,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h10,8'hc,8'h9,8'h10,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'ha,8'h5,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'ha,8'hd,8'hd,8'hd,8'h7,8'h5,8'h5,8'h17,8'hd,8'hd,8'h17,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h10,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'ha,8'h17,8'h13,8'h17,8'h3,8'h5,8'h5,8'h3,8'hd,8'hd,8'h3,8'ha,8'ha,8'h7,8'h7,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h10,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'ha,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'ha,8'h3,8'h17,8'h3,8'h7,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'ha,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'ha,8'h5,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h3,8'h17,8'h17,8'h17,8'h3,8'h3,8'h3,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'ha,8'h17,8'h12,8'h17,8'ha,8'h10,8'h5,8'h3,8'hd,8'h13,8'h17,8'ha,8'h5,8'ha,8'h7,8'h7,8'h7,8'h3,8'h3,8'h17,8'h3,8'h3,8'h3,8'h3,8'h3,8'h17,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'ha,8'h17,8'h12,8'h17,8'h7,8'h5,8'h5,8'h3,8'hd,8'h13,8'h3,8'ha,8'h5,8'h5,8'ha,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'ha,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'h17,8'h3,8'h7,8'h5,8'h5,8'h3,8'h17,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'h3,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h3,8'h3,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'ha,8'ha,8'ha,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'h8,8'h2,8'h2,8'h2,8'h2,8'h8,8'h8,8'h8,8'h8,8'h8,8'ha,8'h3,8'h17,8'h3,8'ha,8'h5,8'h5,8'h3,8'h3,8'h17,8'h3,8'ha,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'ha,8'h17,8'h12,8'h17,8'ha,8'h5,8'h5,8'h3,8'hd,8'h12,8'h17,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'hc,8'h9,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h7,8'h17,8'hd,8'h17,8'h7,8'h5,8'h5,8'h3,8'h17,8'hd,8'h3,8'ha,8'h10,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h5,8'h10,8'h5,8'hc,8'h9,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'hd,8'hd,8'hd,8'hd,8'hd,8'h10,8'h5,8'hd,8'hd,8'hd,8'hd,8'h5,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'h10,8'hc,8'h9};

																																																			                                                                                                                                                                             // Main sprite/////ASH1 = '{ 8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h1,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h1,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h3,8'h3,8'h1,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h1,8'h1,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h3,8'h1,8'h1,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h1,8'h1,8'h1,8'h1,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h3,8'h1,8'h1,8'h1,8'h3,8'h7,8'h7,8'h7,8'h3,8'h2,8'h3,8'h7,8'h7,8'h7,8'h1,8'h1,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h3,8'h1,8'h1,8'h1,8'h3,8'h7,8'h3,8'h3,8'h2,8'h2,8'h3,8'h3,8'h7,8'h7,8'h1,8'h1,8'h1,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h3,8'h1,8'h1,8'h1,8'h3,8'h7,8'h2,8'h3,8'h7,8'h7,8'h7,8'h2,8'h3,8'h7,8'h1,8'h1,8'h1,8'h3,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h1,8'h3,8'h7,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h7,8'h7,8'h1,8'h1,8'h3,8'h3,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h1,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h1,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h1,8'h3,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h3,8'h4,8'h3,8'h3,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h4,8'h4,8'h3,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h3,8'h5,8'h4,8'h4,8'h5,8'h4,8'h7,8'h3,8'h5,8'h5,8'h4,8'h7,8'h4,8'h5,8'h4,8'h4,8'h4,8'h4,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h3,8'h4,8'h4,8'h4,8'h5,8'h4,8'h7,8'h3,8'h5,8'h5,8'h4,8'h7,8'h3,8'h5,8'h4,8'h4,8'h4,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h3,8'h3,8'h4,8'h4,8'h4,8'h3,8'h4,8'h5,8'h5,8'h4,8'h3,8'h4,8'h4,8'h4,8'h4,8'h4,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h3,8'h3,8'h4,8'h1,8'h4,8'h5,8'h5,8'h4,8'h1,8'h4,8'h4,8'h3,8'h3,8'h3,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h1,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h1,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h1,8'h4,8'h3,8'h7,8'h7,8'h7,8'h3,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h4,8'h4,8'h3,8'h0,8'h0,8'h0,8'h0,8'h3,8'h4,8'h5,8'h3,8'h7,8'h7,8'h7,8'h3,8'h6,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h6,8'h6,8'h3,8'h7,8'h7,8'h3,8'h5,8'h4,8'h3,8'h0,8'h0,8'h0,8'h0,8'h3,8'h1,8'h5,8'h4,8'h4,8'h3,8'h7,8'h3,8'h6,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h6,8'h6,8'h3,8'h7,8'h3,8'h4,8'h5,8'h4,8'h3,8'h0,8'h0,8'h0,8'h0,8'h3,8'h1,8'h1,8'h4,8'h4,8'h3,8'h7,8'h3,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h7,8'h7,8'h3,8'h4,8'h4,8'h1,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h6,8'h6,8'h3,8'h1,8'h1,8'h3,8'h6,8'h6,8'h3,8'h3,8'h7,8'h7,8'h7,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h7,8'h7,8'h3,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h0,8'h0,8'h0,8'h3,8'h3,8'h7,8'h7,8'h7,8'h7,8'h3,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h7,8'h7,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h7,8'h7,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0};
																																																			                                                                                                                                                                    			//ASH1 = '{8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h1,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'hf,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h1,8'h16,8'h16,8'h16,8'h16,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h9,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h16,8'h16,8'h1,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h1,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h1,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h16,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'hb,8'hb,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'h11,8'h3,8'h3,8'h3,8'h3,8'h9,8'h11,8'h11,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h11,8'h11,8'h9,8'h3,8'h3,8'h3,8'h3,8'h11,8'hb,8'hb,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'h3,8'hb,8'hb,8'hb,8'hb,8'h9,8'h11,8'h11,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h3,8'h11,8'h11,8'h9,8'h3,8'h3,8'hb,8'hb,8'h3,8'hb,8'hb,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h9,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'h9,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h9,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'h9,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h1,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h1,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h3,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h17,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h3,8'hd,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'hd,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h4,8'h9,8'h4,8'h3,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h7,8'h9,8'h9,8'h4,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'hd,8'h9,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h3,8'h9,8'hd,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h4,8'h4,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h3,8'h11,8'h9,8'hd,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h7,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'hd,8'h3,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h9,8'h9,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'h11,8'h3,8'h11,8'h11,8'h9,8'h9,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h9,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h2,8'h2,8'h11,8'hb,8'hb,8'hb,8'hb,8'h11,8'h11,8'h2,8'h11,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h9,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h9,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h9,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h9,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h9,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h9,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h9,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h9,8'h9,8'h11,8'hf,8'hf,8'h11,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h11,8'hf,8'hf,8'h11,8'h9,8'h9,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hb,8'hb,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'hb,8'hb,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'hb,8'hb,8'hb,8'hb,8'hb,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h7,8'hf,8'hf,8'hf,8'hf,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h11,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hf,8'hf,8'hf,8'hf,8'h11,8'h3,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h11,8'h11,8'h11,8'h11,8'h11,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'hd,8'h11,8'hf,8'hf,8'hf,8'hf,8'hf,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'hf,8'hf,8'hf,8'h11,8'h7,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h11,8'hf,8'hf,8'hf,8'hf,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'hf,8'hf,8'h11,8'h17,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h3,8'h11,8'hf,8'hf,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h17,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h3,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h7,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h11,8'h11,8'h11,8'h11,8'h11,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h11,8'h0,8'h11,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h0,8'h0,8'h0,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h2,8'h2,8'h2,8'h2,8'h2,8'h2,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h2,8'h2,8'h2,8'h2,8'h2,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h16,8'h16,8'h11,8'h11,8'h16,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h16,8'h16,8'h11,8'h11,8'h16,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h16,8'h3,8'h3,8'h16,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h3,8'h16,8'h3,8'h3,8'h16,8'h3,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0,8'h0};

																																																			                                                                                                                                                                    ashDown0 = '{ 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h1, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h15, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h11, 8'h16, 8'h16, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h1, 8'h16, 8'h11, 8'h11, 8'h15, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h11, 8'h16, 8'h1, 8'h3, 8'h11, 8'h11, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'h13, 8'hd, 8'hd, 8'h11, 8'hd, 8'hd, 8'hd, 8'h11, 8'hd, 8'hd, 8'h13, 8'h17, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h13, 8'h13, 8'h14, 8'h14, 8'h3, 8'h14, 8'h14, 8'h14, 8'h3, 8'h14, 8'h14, 8'h13, 8'h13, 8'hd, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h13, 8'h17, 8'h14, 8'h14, 8'h14, 8'h17, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'hd, 8'h13, 8'h13, 8'h17, 8'h14, 8'h14, 8'h14, 8'h17, 8'h13, 8'h13, 8'hd, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h17, 8'h11, 8'h11, 8'h2, 8'h2, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h2, 8'h2, 8'h11, 8'h11, 8'h11, 8'hd, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h14, 8'h13, 8'h17, 8'h11, 8'h2, 8'h2, 8'ha, 8'ha, 8'ha, 8'ha, 8'ha, 8'h2, 8'h2, 8'h11, 8'h17, 8'hd, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h14, 8'h11, 8'h2, 8'h2, 8'h8, 8'h8, 8'h8, 8'h8, 8'h8, 8'h2, 8'h2, 8'h11, 8'h14, 8'h14, 8'h13, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'hd, 8'h11, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h11, 8'hd, 8'hd, 8'h13, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h11, 8'h11, 8'h2, 8'h2, 8'h2, 8'h16, 8'h16, 8'h16, 8'h2, 8'h2, 8'h2, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
																																																			                                                                                                                                                                    ashDown1 = '{ 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h1, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h15, 8'h15, 8'h7, 8'h11, 8'h11, 8'h3, 8'h16, 8'h1, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h15, 8'h15, 8'h7, 8'h11, 8'h11, 8'h3, 8'h16, 8'h1, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h1, 8'h16, 8'h3, 8'h11, 8'h15, 8'h11, 8'h11, 8'h7, 8'h15, 8'h11, 8'h3, 8'h16, 8'h1, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h13, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h13, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h13, 8'h13, 8'h14, 8'h14, 8'h3, 8'h14, 8'h14, 8'h17, 8'h3, 8'h14, 8'h13, 8'h13, 8'hd, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h13, 8'h13, 8'h14, 8'h14, 8'h3, 8'h14, 8'h14, 8'h17, 8'h3, 8'h14, 8'h13, 8'h13, 8'hd, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h13, 8'h13, 8'h17, 8'h14, 8'h14, 8'hd, 8'h17, 8'h13, 8'h13, 8'h13, 8'h17, 8'h11, 8'h17, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h13, 8'h13, 8'h17, 8'h14, 8'h14, 8'hd, 8'h17, 8'h13, 8'h13, 8'h13, 8'h17, 8'h11, 8'h17, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'hd, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h17, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'ha, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'ha, 8'h2, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'ha, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'ha, 8'h2, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h14, 8'h14, 8'hd, 8'h17, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h13, 8'h13, 8'h1, 8'h17, 8'h2, 8'h16, 8'h16, 8'h16, 8'h2, 8'h8, 8'ha, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h13, 8'h13, 8'h1, 8'h17, 8'h2, 8'h16, 8'h16, 8'h16, 8'h2, 8'h8, 8'ha, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
																																																			                                                                                                                                                                    ashDown2 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h16, 8'h16, 8'h11, 8'h11, 8'h7, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h3, 8'h16, 8'h16, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'hd, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h3, 8'h13, 8'h13, 8'h14, 8'hd, 8'h3, 8'h14, 8'h14, 8'h12, 8'h11, 8'h14, 8'h13, 8'h13, 8'h13, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h3, 8'h13, 8'h13, 8'h14, 8'hd, 8'h3, 8'h14, 8'h14, 8'h12, 8'h11, 8'h14, 8'h13, 8'h13, 8'h13, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h17, 8'h11, 8'h17, 8'hd, 8'h13, 8'hd, 8'hd, 8'h14, 8'h14, 8'h14, 8'h17, 8'h13, 8'h13, 8'h1, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h17, 8'h11, 8'h17, 8'hd, 8'h13, 8'hd, 8'hd, 8'h14, 8'h14, 8'h14, 8'h17, 8'h13, 8'h13, 8'h1, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h17, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h2, 8'h8, 8'ha, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h2, 8'h8, 8'ha, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h3, 8'hd, 8'h14, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h2, 8'h2, 8'hd, 8'h16, 8'h16, 8'h16, 8'h2, 8'h17, 8'hd, 8'h13, 8'h13, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h2, 8'h2, 8'hd, 8'h16, 8'h16, 8'h16, 8'h2, 8'h17, 8'hd, 8'h13, 8'h13, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0 };

																																																			                                                                                                                                                                    ashLeft0 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h15, 8'h15, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h1, 8'h1, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h3, 8'h3, 8'h17, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h1, 8'h17, 8'h17, 8'h17, 8'h1, 8'h17, 8'h17, 8'h17, 8'h1, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h11, 8'h13, 8'h13, 8'h13, 8'h17, 8'h14, 8'h13, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h11, 8'h13, 8'h13, 8'h13, 8'h17, 8'h14, 8'h13, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h14, 8'h14, 8'h3, 8'h14, 8'h13, 8'h13, 8'hd, 8'h14, 8'h13, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'hd, 8'h14, 8'h13, 8'h13, 8'h14, 8'h13, 8'hd, 8'hd, 8'h7, 8'h11, 8'h11, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'hd, 8'hd, 8'hd, 8'hd, 8'h17, 8'h3, 8'h17, 8'h17, 8'h15, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h17, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h8, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'ha, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'hd, 8'h7, 8'h7, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h14, 8'h14, 8'h14, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'hd, 8'hd, 8'hd, 8'h11, 8'h11, 8'h11, 8'h7, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h3, 8'h3, 8'h3, 8'h17, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
																																																			                                                                                                                                                                    ashLeft1 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h15, 8'h7, 8'h11, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h15, 8'h7, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h15, 8'h7, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h17, 8'h1, 8'h1, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h3, 8'h3, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h1, 8'h3, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h14, 8'h3, 8'h17, 8'h14, 8'h13, 8'h17, 8'h14, 8'h14, 8'h14, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h17, 8'h14, 8'h17, 8'hd, 8'h14, 8'h13, 8'h13, 8'h14, 8'h14, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'hd, 8'h13, 8'h13, 8'h13, 8'h13, 8'hd, 8'hd, 8'h1, 8'h7, 8'h7, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h17, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'hd, 8'hd, 8'hd, 8'h17, 8'h17, 8'h17, 8'h17, 8'hd, 8'h15, 8'h15, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h17, 8'h17, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h13, 8'h12, 8'h13, 8'h11, 8'h11, 8'h11, 8'h2, 8'h2, 8'h15, 8'h15, 8'h15, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h11, 8'h14, 8'h14, 8'h12, 8'h11, 8'h11, 8'h11, 8'h2, 8'h8, 8'h15, 8'h15, 8'he, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h14, 8'h14, 8'h13, 8'h11, 8'h11, 8'h11, 8'h2, 8'h2, 8'h7, 8'h17, 8'he, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h13, 8'h13, 8'hd, 8'h11, 8'h11, 8'h11, 8'h2, 8'h2, 8'h11, 8'h17, 8'he, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
																																																			                                                                                                                                                                    ashLeft2 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h17, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h1, 8'h15, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h1, 8'h15, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h17, 8'h3, 8'h3, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h1, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h1, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h16, 8'h3, 8'h3, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h3, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h17, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h17, 8'h17, 8'h11, 8'h3, 8'h17, 8'h17, 8'h3, 8'h3, 8'hd, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h14, 8'h11, 8'hd, 8'h14, 8'h14, 8'hd, 8'hd, 8'h14, 8'h13, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h14, 8'h3, 8'hd, 8'h14, 8'h13, 8'h13, 8'h13, 8'h14, 8'h13, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h14, 8'h17, 8'hd, 8'h14, 8'h13, 8'h13, 8'h13, 8'h14, 8'h13, 8'h17, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h15, 8'h15, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h17, 8'h3, 8'h3, 8'h3, 8'h11, 8'he, 8'h15, 8'h15, 8'he, 8'he, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h6, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h3, 8'h12, 8'h15, 8'h15, 8'he, 8'h7, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h2, 8'h2, 8'h8, 8'h11, 8'h11, 8'h3, 8'h14, 8'h14, 8'h12, 8'h15, 8'h17, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'ha, 8'h2, 8'h11, 8'h11, 8'h3, 8'h13, 8'h13, 8'h17, 8'h17, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'ha, 8'h2, 8'h3, 8'h11, 8'h3, 8'hd, 8'h13, 8'hd, 8'h17, 8'h15, 8'h15, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h11, 8'h11, 8'h3, 8'h12, 8'h15, 8'h15, 8'hf, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h7, 8'h7, 8'h7, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};

																																																			                                                                                                                                                                    ashRight0 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h7, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h11, 8'h15, 8'h15, 8'h1, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h7, 8'he, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h1, 8'h1, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'hd, 8'h13, 8'h13, 8'h3, 8'hd, 8'hd, 8'hd, 8'h11, 8'hd, 8'hd, 8'hd, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h14, 8'h14, 8'h17, 8'h13, 8'h13, 8'h13, 8'h11, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h14, 8'h14, 8'h13, 8'h13, 8'h14, 8'h14, 8'h3, 8'h14, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h14, 8'h14, 8'h13, 8'h13, 8'h14, 8'h14, 8'h17, 8'h14, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h17, 8'h17, 8'h1, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'hf, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h2, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h17, 8'he, 8'hd, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h8, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h15, 8'he, 8'h17, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h2, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'h15, 8'h15, 8'h11, 8'h11, 8'h3, 8'h13, 8'h13, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h11, 8'h11, 8'h3, 8'h13, 8'h13, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h17, 8'h17, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0 };
																																																			                                                                                                                                                                    ashRight1 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'hf, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h15, 8'h3, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h15, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h15, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h11, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h1, 8'h16, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'hd, 8'h13, 8'h14, 8'h3, 8'hd, 8'h13, 8'hd, 8'hd, 8'h11, 8'h13, 8'h13, 8'h13, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h13, 8'h13, 8'h14, 8'hd, 8'h13, 8'h13, 8'h14, 8'h14, 8'h3, 8'h14, 8'hd, 8'h1, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'hf, 8'h13, 8'h13, 8'h14, 8'h13, 8'h13, 8'h13, 8'h14, 8'h12, 8'h17, 8'h14, 8'hd, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h17, 8'h11, 8'h15, 8'hd, 8'hd, 8'hd, 8'h13, 8'h13, 8'h13, 8'h14, 8'h13, 8'hd, 8'hd, 8'hd, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hd, 8'h11, 8'h15, 8'h17, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h15, 8'h15, 8'h15, 8'h17, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h15, 8'h15, 8'h15, 8'h17, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h17, 8'h15, 8'h15, 8'h15, 8'ha, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'hd, 8'h17, 8'h17, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h17, 8'he, 8'h7, 8'hd, 8'h8, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h14, 8'h14, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h15, 8'h3, 8'h11, 8'h11, 8'h2, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h13, 8'h13, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'hd, 8'h15, 8'he, 8'h11, 8'h11, 8'h2, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'hd, 8'hd, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h15, 8'h7, 8'h11, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h3, 8'h1, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
																																																			                                                                                                                                                                    ashRight2 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'hf, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h7, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h15, 8'h1, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h15, 8'h1, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h1, 8'h17, 8'h1, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h3, 8'h3, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h3, 8'h1, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h1, 8'h17, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h17, 8'h3, 8'h3, 8'h17, 8'h17, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h13, 8'h14, 8'h17, 8'h17, 8'h14, 8'h14, 8'h11, 8'h11, 8'h14, 8'h14, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h13, 8'h14, 8'h17, 8'h17, 8'h13, 8'h13, 8'h3, 8'h11, 8'h13, 8'h13, 8'hd, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h13, 8'h14, 8'h13, 8'h13, 8'h13, 8'h14, 8'h17, 8'h17, 8'h14, 8'h14, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h15, 8'he, 8'h17, 8'h17, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h13, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h7, 8'h7, 8'h15, 8'h15, 8'he, 8'h11, 8'h3, 8'h3, 8'h3, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h3, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'he, 8'he, 8'h15, 8'h15, 8'h12, 8'h3, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'h15, 8'h12, 8'h14, 8'h14, 8'h11, 8'h11, 8'h11, 8'h2, 8'h2, 8'h2, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h17, 8'he, 8'hd, 8'h14, 8'h14, 8'h11, 8'h11, 8'h11, 8'h2, 8'ha, 8'ha, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h15, 8'h15, 8'h17, 8'h1, 8'h13, 8'h13, 8'h11, 8'h11, 8'h11, 8'h8, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'hf, 8'hf, 8'he, 8'h15, 8'h12, 8'h3, 8'h11, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h7, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};

																																																			                                                                                                                                                                    ashUp0 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h17, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h1, 8'h17, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h17, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h3, 8'h7, 8'h7, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h7, 8'h3, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h17, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h17, 8'h3, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h14, 8'h14, 8'h11, 8'h2, 8'h15, 8'h15, 8'h8, 8'h8, 8'h8, 8'h8, 8'h8, 8'h8, 8'h15, 8'h2, 8'ha, 8'h11, 8'h14, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h14, 8'h14, 8'h11, 8'h2, 8'h15, 8'h15, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'h15, 8'h2, 8'ha, 8'h11, 8'h14, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h17, 8'h8, 8'h17, 8'h17, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h17, 8'h8, 8'ha, 8'h17, 8'h13, 8'h17, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h11, 8'h11, 8'he, 8'he, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'he, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h17, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h3, 8'h3, 8'h15, 8'h3, 8'h3, 8'h3, 8'h15, 8'h15, 8'h3, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
																																																			                                                                                                                                                                    ashUp1 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h1, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h1, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h17, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h3, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h1, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h17, 8'h1, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h1, 8'h1, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h17, 8'h3, 8'h11, 8'h11, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h17, 8'h17, 8'h15, 8'h2, 8'h8, 8'h8, 8'h8, 8'h8, 8'h8, 8'h15, 8'h2, 8'h2, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'hd, 8'h17, 8'h11, 8'h2, 8'h2, 8'h17, 8'h5, 8'h5, 8'h5, 8'h5, 8'h5, 8'h5, 8'h17, 8'h2, 8'h2, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h13, 8'hd, 8'h11, 8'h2, 8'h2, 8'h17, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h3, 8'h2, 8'h2, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h13, 8'h13, 8'h13, 8'h8, 8'h2, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h2, 8'h8, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'hf, 8'h15, 8'h15, 8'hd, 8'hd, 8'h15, 8'h15, 8'hf, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h7, 8'h7, 8'h3, 8'h3, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h1, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
																																																			                                                                                                                                                                    ashUp2 = '{8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h17, 8'h17, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h17, 8'h3, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h7, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h7, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h16, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h1, 8'h1, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h1, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h16, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h16, 8'h16, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h13, 8'h13, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h17, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h17, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h11, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h17, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h2, 8'h15, 8'hd, 8'h2, 8'h2, 8'h2, 8'h2, 8'h2, 8'hd, 8'h15, 8'h3, 8'h3, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h2, 8'he, 8'hd, 8'h5, 8'h5, 8'h5, 8'h5, 8'h5, 8'hd, 8'h17, 8'h2, 8'h2, 8'h11, 8'h17, 8'hd, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h17, 8'h17, 8'h2, 8'h3, 8'h17, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h17, 8'h3, 8'h2, 8'h2, 8'h11, 8'h13, 8'h13, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h8, 8'he, 8'he, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'he, 8'he, 8'h8, 8'h8, 8'h17, 8'h13, 8'h13, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'ha, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'ha, 8'ha, 8'hd, 8'h1, 8'hd, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h11, 8'h11, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h3, 8'h11, 8'h15, 8'h15, 8'h15, 8'he, 8'h15, 8'he, 8'h15, 8'h15, 8'h15, 8'h11, 8'h11, 8'h3, 8'h3, 8'h17, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h7, 8'h15, 8'h17, 8'h17, 8'h17, 8'h15, 8'h7, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h3, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h1, 8'h17, 8'h17, 8'h11, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h3, 8'h11, 8'h11, 8'h11, 8'h3, 8'h3, 8'h3, 8'h3, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h11, 8'h11, 8'h11, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0};
																																																			                                                                                                                                                                    				 end



																																																			                                                                                                                                                                    */

//colorTable c0();

//spriteTable s0();

// Compute whether the pixel corresponds to ball or background\


//////////////////Uncomment from here//////////////////
//always_comb
//begin : Ball_on_proc
//if ( ( DistX >= 0 && DistX <= 28  && DistY >= 0 && DistY <= 40))
//       ash_on= 1'b1;
//              else
//              ash_on = 1'b0;
//end
//
//// Assign color based on ball_on signal
//always_comb
//begin : RGB_Display
//if ((ash_on == 1'b1) && ashDown0[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b00 && counter[3:2] == 2'b00  )
//        begin
//        color = ashDown0[DistY*28 +DistX];
//        end
//
//else if ((ash_on == 1'b1) && ashDown1[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b00 && counter[3:2] == 2'b01 )
//        begin
//        color = ashDown1[DistY*28 +DistX];
//        end
//
//else if ((ash_on == 1'b1) && ashDown2[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b00 && counter[3:2] == 2'b10 )
//        begin
//        color = ashDown2[DistY*28 +DistX];
//        end
//
//else if ((ash_on == 1'b1) && ashLeft0[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b01 && counter[3:2] == 2'b00 )
//        begin
//        color = ashLeft0[DistY*28 +DistX];
//        end
//
//else if ((ash_on == 1'b1) && ashLeft1[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b01 && counter[3:2] == 2'b01)
//        begin
//        color = ashLeft1[DistY*28 +DistX];
//        end
//
//else if ((ash_on == 1'b1) && ashLeft2[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b01 && counter[3:2] == 2'b10)
//        begin
//        color = ashLeft2[DistY*28 +DistX];
//        end
//
//else if ((ash_on == 1'b1) && ashRight0[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b10 && counter[3:2] == 2'b00 )
//        begin
//        color = ashRight0[DistY*28 +DistX];
//        end
//
//else if ((ash_on == 1'b1) && ashRight1[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b10 && counter[3:2] == 2'b01)
//        begin
//        color = ashRight1[DistY*28 +DistX];
//        end
//
//else if ((ash_on == 1'b1) && ashRight2[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b10 && counter[3:2] == 2'b10)
//        begin
//        color = ashRight2[DistY*28 +DistX];
//        end
//
//else if ((ash_on == 1'b1) && ashUp0[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b11 && counter[3:2] == 2'b00 )
//        begin
//        color = ashUp0[DistY*28 +DistX];
//        end
//
//else if ((ash_on == 1'b1) && ashUp1[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b11 && counter[3:2] == 2'b01)
//        begin
//        color = ashUp1[DistY*28 +DistX];
//        end
//
//else if ((ash_on == 1'b1) && ashUp2[DistY*28 +DistX]!=8'h0 && spriteDirControl == 2'b11 && counter[3:2] == 2'b10)
//        begin
//        color = ashUp2[DistY*28 +DistX];
//        end
//
//        else
//            begin
//				//color = color[pixel];
//				//color = MAP1[pixel];
//				color = Data;
//				end
//        end

//////////////////Uncomment from here//////////////////

																																																			                                                                                                                                                                    //else if( DrawX >= 42 && DrawX <= 146 && DrawY == 66 ) // Poke center top border
//		  begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawX >=42 && DrawX<=146 && DrawY== 146) //Poke center bottom border
//		  begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawY >=66 && DrawY<=146 && DrawX== 42) //Poke center left border
//		  begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawY >=66 && DrawY<=146 && DrawX== 146) //Poke center right border
//		  begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawX==0 && DrawY==30) // Left top corner of the map
//         begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawX==10 && DrawY==30) // Left top corner of the map
//         begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawX==20 && DrawY==30) // Left top corner of the map
//         begin
//		  color = 8'd0;
//		  end
//
//		  else if(DrawX==30 && DrawY==30) // Left top corner of the map
//         begin
//		  color = 8'd0;
//		  end
//
//		   else if(DrawX==0 && DrawY==480)    //Left bottom corner of the map
//         begin
//		  color = 8'd0;
//		  end
//
//		   else if(DrawX==640 && DrawY==0) // Right top corner
//         begin
//		  color = 8'd0;
//		  end
//
//		   else if(DrawX==640 && DrawY==480) // Right bottom
//         begin
//		  color = 8'd0;
//		  end
//
//int pixel;




//        endmodule


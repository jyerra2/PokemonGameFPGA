module starterSelect(input logic [1:0] starterSelect,
							input logic [4:0] prev_ID,
							input logic enable,
							output logic [4:0] new_ID); 